VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32_1RW1R
  CLASS BLOCK ;
  FOREIGN RAM32_1RW1R ;
  ORIGIN 0.000 0.000 ;
  SIZE 1274.560 BY 160.720 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 87.920 1274.560 88.480 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 103.600 1274.560 104.160 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 119.280 1274.560 119.840 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 134.960 1274.560 135.520 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 150.640 1274.560 151.200 ;
    END
  END A0[4]
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.160 2.000 34.720 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 2.000 57.680 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.080 2.000 80.640 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.040 2.000 103.600 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 2.000 126.560 ;
    END
  END A1[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.200 2.000 11.760 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.720 0.000 21.280 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.320 0.000 418.880 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 0.000 458.640 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.840 0.000 498.400 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.360 0.000 577.920 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 0.000 617.680 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 656.880 0.000 657.440 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 736.400 0.000 736.960 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 815.920 0.000 816.480 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 855.680 0.000 856.240 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 895.440 0.000 896.000 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 0.000 935.760 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.960 0.000 975.520 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 0.000 1015.280 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1054.480 0.000 1055.040 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1094.240 0.000 1094.800 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1134.000 0.000 1134.560 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1173.760 0.000 1174.320 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.240 0.000 100.800 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1213.520 0.000 1214.080 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1253.280 0.000 1253.840 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.760 0.000 180.320 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.280 0.000 259.840 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 0.000 339.360 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.600 158.720 20.160 160.720 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 158.720 216.160 160.720 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 158.720 255.360 160.720 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.000 158.720 294.560 160.720 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.200 158.720 333.760 160.720 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 158.720 372.960 160.720 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.600 158.720 412.160 160.720 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.800 158.720 451.360 160.720 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.000 158.720 490.560 160.720 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.200 158.720 529.760 160.720 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.400 158.720 568.960 160.720 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 158.720 39.760 160.720 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.600 158.720 608.160 160.720 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 627.200 158.720 627.760 160.720 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.800 158.720 647.360 160.720 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 158.720 666.960 160.720 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.000 158.720 686.560 160.720 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 158.720 706.160 160.720 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.200 158.720 725.760 160.720 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.800 158.720 745.360 160.720 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 764.400 158.720 764.960 160.720 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 784.000 158.720 784.560 160.720 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 158.720 59.360 160.720 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.600 158.720 804.160 160.720 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 158.720 823.760 160.720 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 158.720 78.960 160.720 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 158.720 98.560 160.720 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 158.720 118.160 160.720 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.200 158.720 137.760 160.720 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 158.720 157.360 160.720 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.400 158.720 176.960 160.720 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 158.720 196.560 160.720 ;
    END
  END Do0[9]
  PIN Do1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 158.720 235.760 160.720 ;
    END
  END Do1[0]
  PIN Do1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 842.800 158.720 843.360 160.720 ;
    END
  END Do1[10]
  PIN Do1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 158.720 862.960 160.720 ;
    END
  END Do1[11]
  PIN Do1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 882.000 158.720 882.560 160.720 ;
    END
  END Do1[12]
  PIN Do1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 158.720 902.160 160.720 ;
    END
  END Do1[13]
  PIN Do1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 921.200 158.720 921.760 160.720 ;
    END
  END Do1[14]
  PIN Do1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 158.720 941.360 160.720 ;
    END
  END Do1[15]
  PIN Do1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.400 158.720 960.960 160.720 ;
    END
  END Do1[16]
  PIN Do1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 980.000 158.720 980.560 160.720 ;
    END
  END Do1[17]
  PIN Do1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 999.600 158.720 1000.160 160.720 ;
    END
  END Do1[18]
  PIN Do1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 158.720 1019.760 160.720 ;
    END
  END Do1[19]
  PIN Do1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 158.720 274.960 160.720 ;
    END
  END Do1[1]
  PIN Do1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1038.800 158.720 1039.360 160.720 ;
    END
  END Do1[20]
  PIN Do1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 158.720 1058.960 160.720 ;
    END
  END Do1[21]
  PIN Do1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1078.000 158.720 1078.560 160.720 ;
    END
  END Do1[22]
  PIN Do1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1097.600 158.720 1098.160 160.720 ;
    END
  END Do1[23]
  PIN Do1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1117.200 158.720 1117.760 160.720 ;
    END
  END Do1[24]
  PIN Do1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1136.800 158.720 1137.360 160.720 ;
    END
  END Do1[25]
  PIN Do1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1156.400 158.720 1156.960 160.720 ;
    END
  END Do1[26]
  PIN Do1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1176.000 158.720 1176.560 160.720 ;
    END
  END Do1[27]
  PIN Do1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1195.600 158.720 1196.160 160.720 ;
    END
  END Do1[28]
  PIN Do1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1215.200 158.720 1215.760 160.720 ;
    END
  END Do1[29]
  PIN Do1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 158.720 314.160 160.720 ;
    END
  END Do1[2]
  PIN Do1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1234.800 158.720 1235.360 160.720 ;
    END
  END Do1[30]
  PIN Do1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1254.400 158.720 1254.960 160.720 ;
    END
  END Do1[31]
  PIN Do1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 158.720 353.360 160.720 ;
    END
  END Do1[3]
  PIN Do1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 158.720 392.560 160.720 ;
    END
  END Do1[4]
  PIN Do1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 158.720 431.760 160.720 ;
    END
  END Do1[5]
  PIN Do1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 158.720 470.960 160.720 ;
    END
  END Do1[6]
  PIN Do1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 158.720 510.160 160.720 ;
    END
  END Do1[7]
  PIN Do1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 158.720 549.360 160.720 ;
    END
  END Do1[8]
  PIN Do1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 158.720 588.560 160.720 ;
    END
  END Do1[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 9.520 1274.560 10.080 ;
    END
  END EN0
  PIN EN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 2.000 149.520 ;
    END
  END EN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 18.320 11.460 19.920 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 171.920 11.460 173.520 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 325.520 11.460 327.120 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 479.120 11.460 480.720 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 632.720 11.460 634.320 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 786.320 11.460 787.920 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 939.920 11.460 941.520 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1093.520 11.460 1095.120 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1247.120 11.460 1248.720 149.260 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 95.120 11.460 96.720 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 248.720 11.460 250.320 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 402.320 11.460 403.920 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.920 11.460 557.520 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 709.520 11.460 711.120 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 863.120 11.460 864.720 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1016.720 11.460 1018.320 149.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1170.320 11.460 1171.920 149.260 ;
    END
  END VSS
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 25.200 1274.560 25.760 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 40.880 1274.560 41.440 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 56.560 1274.560 57.120 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1272.560 72.240 1274.560 72.800 ;
    END
  END WE0[3]
  OBS
      LAYER Metal1 ;
        RECT 2.330 0.150 1271.760 160.570 ;
      LAYER Metal2 ;
        RECT 0.140 158.420 19.300 160.630 ;
        RECT 20.460 158.420 38.900 160.630 ;
        RECT 40.060 158.420 58.500 160.630 ;
        RECT 59.660 158.420 78.100 160.630 ;
        RECT 79.260 158.420 97.700 160.630 ;
        RECT 98.860 158.420 117.300 160.630 ;
        RECT 118.460 158.420 136.900 160.630 ;
        RECT 138.060 158.420 156.500 160.630 ;
        RECT 157.660 158.420 176.100 160.630 ;
        RECT 177.260 158.420 195.700 160.630 ;
        RECT 196.860 158.420 215.300 160.630 ;
        RECT 216.460 158.420 234.900 160.630 ;
        RECT 236.060 158.420 254.500 160.630 ;
        RECT 255.660 158.420 274.100 160.630 ;
        RECT 275.260 158.420 293.700 160.630 ;
        RECT 294.860 158.420 313.300 160.630 ;
        RECT 314.460 158.420 332.900 160.630 ;
        RECT 334.060 158.420 352.500 160.630 ;
        RECT 353.660 158.420 372.100 160.630 ;
        RECT 373.260 158.420 391.700 160.630 ;
        RECT 392.860 158.420 411.300 160.630 ;
        RECT 412.460 158.420 430.900 160.630 ;
        RECT 432.060 158.420 450.500 160.630 ;
        RECT 451.660 158.420 470.100 160.630 ;
        RECT 471.260 158.420 489.700 160.630 ;
        RECT 490.860 158.420 509.300 160.630 ;
        RECT 510.460 158.420 528.900 160.630 ;
        RECT 530.060 158.420 548.500 160.630 ;
        RECT 549.660 158.420 568.100 160.630 ;
        RECT 569.260 158.420 587.700 160.630 ;
        RECT 588.860 158.420 607.300 160.630 ;
        RECT 608.460 158.420 626.900 160.630 ;
        RECT 628.060 158.420 646.500 160.630 ;
        RECT 647.660 158.420 666.100 160.630 ;
        RECT 667.260 158.420 685.700 160.630 ;
        RECT 686.860 158.420 705.300 160.630 ;
        RECT 706.460 158.420 724.900 160.630 ;
        RECT 726.060 158.420 744.500 160.630 ;
        RECT 745.660 158.420 764.100 160.630 ;
        RECT 765.260 158.420 783.700 160.630 ;
        RECT 784.860 158.420 803.300 160.630 ;
        RECT 804.460 158.420 822.900 160.630 ;
        RECT 824.060 158.420 842.500 160.630 ;
        RECT 843.660 158.420 862.100 160.630 ;
        RECT 863.260 158.420 881.700 160.630 ;
        RECT 882.860 158.420 901.300 160.630 ;
        RECT 902.460 158.420 920.900 160.630 ;
        RECT 922.060 158.420 940.500 160.630 ;
        RECT 941.660 158.420 960.100 160.630 ;
        RECT 961.260 158.420 979.700 160.630 ;
        RECT 980.860 158.420 999.300 160.630 ;
        RECT 1000.460 158.420 1018.900 160.630 ;
        RECT 1020.060 158.420 1038.500 160.630 ;
        RECT 1039.660 158.420 1058.100 160.630 ;
        RECT 1059.260 158.420 1077.700 160.630 ;
        RECT 1078.860 158.420 1097.300 160.630 ;
        RECT 1098.460 158.420 1116.900 160.630 ;
        RECT 1118.060 158.420 1136.500 160.630 ;
        RECT 1137.660 158.420 1156.100 160.630 ;
        RECT 1157.260 158.420 1175.700 160.630 ;
        RECT 1176.860 158.420 1195.300 160.630 ;
        RECT 1196.460 158.420 1214.900 160.630 ;
        RECT 1216.060 158.420 1234.500 160.630 ;
        RECT 1235.660 158.420 1254.100 160.630 ;
        RECT 1255.260 158.420 1273.300 160.630 ;
        RECT 0.140 2.300 1273.300 158.420 ;
        RECT 0.140 0.090 20.420 2.300 ;
        RECT 21.580 0.090 60.180 2.300 ;
        RECT 61.340 0.090 99.940 2.300 ;
        RECT 101.100 0.090 139.700 2.300 ;
        RECT 140.860 0.090 179.460 2.300 ;
        RECT 180.620 0.090 219.220 2.300 ;
        RECT 220.380 0.090 258.980 2.300 ;
        RECT 260.140 0.090 298.740 2.300 ;
        RECT 299.900 0.090 338.500 2.300 ;
        RECT 339.660 0.090 378.260 2.300 ;
        RECT 379.420 0.090 418.020 2.300 ;
        RECT 419.180 0.090 457.780 2.300 ;
        RECT 458.940 0.090 497.540 2.300 ;
        RECT 498.700 0.090 537.300 2.300 ;
        RECT 538.460 0.090 577.060 2.300 ;
        RECT 578.220 0.090 616.820 2.300 ;
        RECT 617.980 0.090 656.580 2.300 ;
        RECT 657.740 0.090 696.340 2.300 ;
        RECT 697.500 0.090 736.100 2.300 ;
        RECT 737.260 0.090 775.860 2.300 ;
        RECT 777.020 0.090 815.620 2.300 ;
        RECT 816.780 0.090 855.380 2.300 ;
        RECT 856.540 0.090 895.140 2.300 ;
        RECT 896.300 0.090 934.900 2.300 ;
        RECT 936.060 0.090 974.660 2.300 ;
        RECT 975.820 0.090 1014.420 2.300 ;
        RECT 1015.580 0.090 1054.180 2.300 ;
        RECT 1055.340 0.090 1093.940 2.300 ;
        RECT 1095.100 0.090 1133.700 2.300 ;
        RECT 1134.860 0.090 1173.460 2.300 ;
        RECT 1174.620 0.090 1213.220 2.300 ;
        RECT 1214.380 0.090 1252.980 2.300 ;
        RECT 1254.140 0.090 1273.300 2.300 ;
      LAYER Metal3 ;
        RECT 1.770 151.500 1273.350 160.580 ;
        RECT 1.770 150.340 1272.260 151.500 ;
        RECT 1.770 149.820 1273.350 150.340 ;
        RECT 2.300 148.660 1273.350 149.820 ;
        RECT 1.770 135.820 1273.350 148.660 ;
        RECT 1.770 134.660 1272.260 135.820 ;
        RECT 1.770 126.860 1273.350 134.660 ;
        RECT 2.300 125.700 1273.350 126.860 ;
        RECT 1.770 120.140 1273.350 125.700 ;
        RECT 1.770 118.980 1272.260 120.140 ;
        RECT 1.770 104.460 1273.350 118.980 ;
        RECT 1.770 103.900 1272.260 104.460 ;
        RECT 2.300 103.300 1272.260 103.900 ;
        RECT 2.300 102.740 1273.350 103.300 ;
        RECT 1.770 88.780 1273.350 102.740 ;
        RECT 1.770 87.620 1272.260 88.780 ;
        RECT 1.770 80.940 1273.350 87.620 ;
        RECT 2.300 79.780 1273.350 80.940 ;
        RECT 1.770 73.100 1273.350 79.780 ;
        RECT 1.770 71.940 1272.260 73.100 ;
        RECT 1.770 57.980 1273.350 71.940 ;
        RECT 2.300 57.420 1273.350 57.980 ;
        RECT 2.300 56.820 1272.260 57.420 ;
        RECT 1.770 56.260 1272.260 56.820 ;
        RECT 1.770 41.740 1273.350 56.260 ;
        RECT 1.770 40.580 1272.260 41.740 ;
        RECT 1.770 35.020 1273.350 40.580 ;
        RECT 2.300 33.860 1273.350 35.020 ;
        RECT 1.770 26.060 1273.350 33.860 ;
        RECT 1.770 24.900 1272.260 26.060 ;
        RECT 1.770 12.060 1273.350 24.900 ;
        RECT 2.300 10.900 1273.350 12.060 ;
        RECT 1.770 10.380 1273.350 10.900 ;
        RECT 1.770 9.220 1272.260 10.380 ;
        RECT 1.770 0.140 1273.350 9.220 ;
      LAYER Metal4 ;
        RECT 3.500 149.560 1103.620 160.630 ;
        RECT 3.500 11.160 18.020 149.560 ;
        RECT 20.220 11.160 94.820 149.560 ;
        RECT 97.020 11.160 171.620 149.560 ;
        RECT 173.820 11.160 248.420 149.560 ;
        RECT 250.620 11.160 325.220 149.560 ;
        RECT 327.420 11.160 402.020 149.560 ;
        RECT 404.220 11.160 478.820 149.560 ;
        RECT 481.020 11.160 555.620 149.560 ;
        RECT 557.820 11.160 632.420 149.560 ;
        RECT 634.620 11.160 709.220 149.560 ;
        RECT 711.420 11.160 786.020 149.560 ;
        RECT 788.220 11.160 862.820 149.560 ;
        RECT 865.020 11.160 939.620 149.560 ;
        RECT 941.820 11.160 1016.420 149.560 ;
        RECT 1018.620 11.160 1093.220 149.560 ;
        RECT 1095.420 11.160 1103.620 149.560 ;
        RECT 3.500 0.090 1103.620 11.160 ;
  END
END RAM32_1RW1R
END LIBRARY

