module RAM32_1RW1R (CLK,
    EN0,
    EN1,
    VDD,
    VSS,
    A0,
    A1,
    Di0,
    Do0,
    Do1,
    WE0);
 input CLK;
 input EN0;
 input EN1;
 input VDD;
 input VSS;
 input [4:0] A0;
 input [4:0] A1;
 input [31:0] Di0;
 output [31:0] Do0;
 output [31:0] Do1;
 input [3:0] WE0;

 wire \A0BUF[0].X ;
 wire \A0BUF[1].X ;
 wire \A0BUF[2].X ;
 wire \A0BUF[3].X ;
 wire \A0BUF[4].X ;
 wire \A1BUF[0].X ;
 wire \A1BUF[1].X ;
 wire \A1BUF[2].X ;
 wire \A1BUF[3].X ;
 wire \A1BUF[4].X ;
 wire \BYTE[0].FLOATBUF0[0].A ;
 wire \BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BYTE[0].FLOATBUF0[0].TE_BN ;
 wire \BYTE[0].FLOATBUF0[0].Z ;
 wire \BYTE[0].FLOATBUF0[1].TE_BN ;
 wire \BYTE[0].FLOATBUF0[1].Z ;
 wire \BYTE[0].FLOATBUF0[2].TE_BN ;
 wire \BYTE[0].FLOATBUF0[2].Z ;
 wire \BYTE[0].FLOATBUF0[3].TE_BN ;
 wire \BYTE[0].FLOATBUF0[3].Z ;
 wire \BYTE[0].FLOATBUF0[4].TE_BN ;
 wire \BYTE[0].FLOATBUF0[4].Z ;
 wire \BYTE[0].FLOATBUF0[5].TE_BN ;
 wire \BYTE[0].FLOATBUF0[5].Z ;
 wire \BYTE[0].FLOATBUF0[6].TE_BN ;
 wire \BYTE[0].FLOATBUF0[6].Z ;
 wire \BYTE[0].FLOATBUF0[7].TE_BN ;
 wire \BYTE[0].FLOATBUF0[7].Z ;
 wire \BYTE[0].FLOATBUF1[0].A ;
 wire \BYTE[0].FLOATBUF1[0].TE_B ;
 wire \BYTE[0].FLOATBUF1[0].TE_BN ;
 wire \BYTE[0].FLOATBUF1[0].Z ;
 wire \BYTE[0].FLOATBUF1[1].TE_BN ;
 wire \BYTE[0].FLOATBUF1[1].Z ;
 wire \BYTE[0].FLOATBUF1[2].TE_BN ;
 wire \BYTE[0].FLOATBUF1[2].Z ;
 wire \BYTE[0].FLOATBUF1[3].TE_BN ;
 wire \BYTE[0].FLOATBUF1[3].Z ;
 wire \BYTE[0].FLOATBUF1[4].TE_BN ;
 wire \BYTE[0].FLOATBUF1[4].Z ;
 wire \BYTE[0].FLOATBUF1[5].TE_BN ;
 wire \BYTE[0].FLOATBUF1[5].Z ;
 wire \BYTE[0].FLOATBUF1[6].TE_BN ;
 wire \BYTE[0].FLOATBUF1[6].Z ;
 wire \BYTE[0].FLOATBUF1[7].TE_BN ;
 wire \BYTE[0].FLOATBUF1[7].Z ;
 wire \BYTE[1].FLOATBUF0[10].A ;
 wire \BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BYTE[1].FLOATBUF0[10].TE_BN ;
 wire \BYTE[1].FLOATBUF0[10].Z ;
 wire \BYTE[1].FLOATBUF0[11].TE_BN ;
 wire \BYTE[1].FLOATBUF0[11].Z ;
 wire \BYTE[1].FLOATBUF0[12].TE_BN ;
 wire \BYTE[1].FLOATBUF0[12].Z ;
 wire \BYTE[1].FLOATBUF0[13].TE_BN ;
 wire \BYTE[1].FLOATBUF0[13].Z ;
 wire \BYTE[1].FLOATBUF0[14].TE_BN ;
 wire \BYTE[1].FLOATBUF0[14].Z ;
 wire \BYTE[1].FLOATBUF0[15].TE_BN ;
 wire \BYTE[1].FLOATBUF0[15].Z ;
 wire \BYTE[1].FLOATBUF0[8].TE_BN ;
 wire \BYTE[1].FLOATBUF0[8].Z ;
 wire \BYTE[1].FLOATBUF0[9].TE_BN ;
 wire \BYTE[1].FLOATBUF0[9].Z ;
 wire \BYTE[1].FLOATBUF1[10].A ;
 wire \BYTE[1].FLOATBUF1[10].TE_B ;
 wire \BYTE[1].FLOATBUF1[10].TE_BN ;
 wire \BYTE[1].FLOATBUF1[10].Z ;
 wire \BYTE[1].FLOATBUF1[11].TE_BN ;
 wire \BYTE[1].FLOATBUF1[11].Z ;
 wire \BYTE[1].FLOATBUF1[12].TE_BN ;
 wire \BYTE[1].FLOATBUF1[12].Z ;
 wire \BYTE[1].FLOATBUF1[13].TE_BN ;
 wire \BYTE[1].FLOATBUF1[13].Z ;
 wire \BYTE[1].FLOATBUF1[14].TE_BN ;
 wire \BYTE[1].FLOATBUF1[14].Z ;
 wire \BYTE[1].FLOATBUF1[15].TE_BN ;
 wire \BYTE[1].FLOATBUF1[15].Z ;
 wire \BYTE[1].FLOATBUF1[8].TE_BN ;
 wire \BYTE[1].FLOATBUF1[8].Z ;
 wire \BYTE[1].FLOATBUF1[9].TE_BN ;
 wire \BYTE[1].FLOATBUF1[9].Z ;
 wire \BYTE[2].FLOATBUF0[16].A ;
 wire \BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BYTE[2].FLOATBUF0[16].TE_BN ;
 wire \BYTE[2].FLOATBUF0[16].Z ;
 wire \BYTE[2].FLOATBUF0[17].TE_BN ;
 wire \BYTE[2].FLOATBUF0[17].Z ;
 wire \BYTE[2].FLOATBUF0[18].TE_BN ;
 wire \BYTE[2].FLOATBUF0[18].Z ;
 wire \BYTE[2].FLOATBUF0[19].TE_BN ;
 wire \BYTE[2].FLOATBUF0[19].Z ;
 wire \BYTE[2].FLOATBUF0[20].TE_BN ;
 wire \BYTE[2].FLOATBUF0[20].Z ;
 wire \BYTE[2].FLOATBUF0[21].TE_BN ;
 wire \BYTE[2].FLOATBUF0[21].Z ;
 wire \BYTE[2].FLOATBUF0[22].TE_BN ;
 wire \BYTE[2].FLOATBUF0[22].Z ;
 wire \BYTE[2].FLOATBUF0[23].TE_BN ;
 wire \BYTE[2].FLOATBUF0[23].Z ;
 wire \BYTE[2].FLOATBUF1[16].A ;
 wire \BYTE[2].FLOATBUF1[16].TE_B ;
 wire \BYTE[2].FLOATBUF1[16].TE_BN ;
 wire \BYTE[2].FLOATBUF1[16].Z ;
 wire \BYTE[2].FLOATBUF1[17].TE_BN ;
 wire \BYTE[2].FLOATBUF1[17].Z ;
 wire \BYTE[2].FLOATBUF1[18].TE_BN ;
 wire \BYTE[2].FLOATBUF1[18].Z ;
 wire \BYTE[2].FLOATBUF1[19].TE_BN ;
 wire \BYTE[2].FLOATBUF1[19].Z ;
 wire \BYTE[2].FLOATBUF1[20].TE_BN ;
 wire \BYTE[2].FLOATBUF1[20].Z ;
 wire \BYTE[2].FLOATBUF1[21].TE_BN ;
 wire \BYTE[2].FLOATBUF1[21].Z ;
 wire \BYTE[2].FLOATBUF1[22].TE_BN ;
 wire \BYTE[2].FLOATBUF1[22].Z ;
 wire \BYTE[2].FLOATBUF1[23].TE_BN ;
 wire \BYTE[2].FLOATBUF1[23].Z ;
 wire \BYTE[3].FLOATBUF0[24].A ;
 wire \BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BYTE[3].FLOATBUF0[24].TE_BN ;
 wire \BYTE[3].FLOATBUF0[24].Z ;
 wire \BYTE[3].FLOATBUF0[25].TE_BN ;
 wire \BYTE[3].FLOATBUF0[25].Z ;
 wire \BYTE[3].FLOATBUF0[26].TE_BN ;
 wire \BYTE[3].FLOATBUF0[26].Z ;
 wire \BYTE[3].FLOATBUF0[27].TE_BN ;
 wire \BYTE[3].FLOATBUF0[27].Z ;
 wire \BYTE[3].FLOATBUF0[28].TE_BN ;
 wire \BYTE[3].FLOATBUF0[28].Z ;
 wire \BYTE[3].FLOATBUF0[29].TE_BN ;
 wire \BYTE[3].FLOATBUF0[29].Z ;
 wire \BYTE[3].FLOATBUF0[30].TE_BN ;
 wire \BYTE[3].FLOATBUF0[30].Z ;
 wire \BYTE[3].FLOATBUF0[31].TE_BN ;
 wire \BYTE[3].FLOATBUF0[31].Z ;
 wire \BYTE[3].FLOATBUF1[24].A ;
 wire \BYTE[3].FLOATBUF1[24].TE_B ;
 wire \BYTE[3].FLOATBUF1[24].TE_BN ;
 wire \BYTE[3].FLOATBUF1[24].Z ;
 wire \BYTE[3].FLOATBUF1[25].TE_BN ;
 wire \BYTE[3].FLOATBUF1[25].Z ;
 wire \BYTE[3].FLOATBUF1[26].TE_BN ;
 wire \BYTE[3].FLOATBUF1[26].Z ;
 wire \BYTE[3].FLOATBUF1[27].TE_BN ;
 wire \BYTE[3].FLOATBUF1[27].Z ;
 wire \BYTE[3].FLOATBUF1[28].TE_BN ;
 wire \BYTE[3].FLOATBUF1[28].Z ;
 wire \BYTE[3].FLOATBUF1[29].TE_BN ;
 wire \BYTE[3].FLOATBUF1[29].Z ;
 wire \BYTE[3].FLOATBUF1[30].TE_BN ;
 wire \BYTE[3].FLOATBUF1[30].Z ;
 wire \BYTE[3].FLOATBUF1[31].TE_BN ;
 wire \BYTE[3].FLOATBUF1[31].Z ;
 wire \CLKBUF.X ;
 wire \DEC0.A_N[0] ;
 wire \DEC0.A_N[1] ;
 wire \DEC0.EN ;
 wire \DEC0.EN_N ;
 wire \DEC1.A_N[0] ;
 wire \DEC1.A_N[1] ;
 wire \DEC1.EN ;
 wire \DEC1.EN_N ;
 wire \DIBUF[0].X ;
 wire \DIBUF[10].X ;
 wire \DIBUF[11].X ;
 wire \DIBUF[12].X ;
 wire \DIBUF[13].X ;
 wire \DIBUF[14].X ;
 wire \DIBUF[15].X ;
 wire \DIBUF[16].X ;
 wire \DIBUF[17].X ;
 wire \DIBUF[18].X ;
 wire \DIBUF[19].X ;
 wire \DIBUF[1].X ;
 wire \DIBUF[20].X ;
 wire \DIBUF[21].X ;
 wire \DIBUF[22].X ;
 wire \DIBUF[23].X ;
 wire \DIBUF[24].X ;
 wire \DIBUF[25].X ;
 wire \DIBUF[26].X ;
 wire \DIBUF[27].X ;
 wire \DIBUF[28].X ;
 wire \DIBUF[29].X ;
 wire \DIBUF[2].X ;
 wire \DIBUF[30].X ;
 wire \DIBUF[31].X ;
 wire \DIBUF[3].X ;
 wire \DIBUF[4].X ;
 wire \DIBUF[5].X ;
 wire \DIBUF[6].X ;
 wire \DIBUF[7].X ;
 wire \DIBUF[8].X ;
 wire \DIBUF[9].X ;
 wire \Do0_REG.CLKBUF[0] ;
 wire \Do0_REG.CLKBUF[1] ;
 wire \Do0_REG.CLKBUF[2] ;
 wire \Do0_REG.CLKBUF[3] ;
 wire \Do0_REG.CLK_buf ;
 wire \Do1_REG.CLKBUF[0] ;
 wire \Do1_REG.CLKBUF[1] ;
 wire \Do1_REG.CLKBUF[2] ;
 wire \Do1_REG.CLKBUF[3] ;
 wire \Do1_REG.CLK_buf ;
 wire \SLICE[0].RAM8.CLKBUF.X ;
 wire \SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[0].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[0].RAM8.DEC0.EN ;
 wire \SLICE[0].RAM8.DEC0.EN_buf ;
 wire \SLICE[0].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[0].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[0].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[0].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[0].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[0].RAM8.DEC1.EN ;
 wire \SLICE[0].RAM8.DEC1.EN_buf ;
 wire \SLICE[0].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[0].RAM8.WEBUF[0].A ;
 wire \SLICE[0].RAM8.WEBUF[0].X ;
 wire \SLICE[0].RAM8.WEBUF[1].A ;
 wire \SLICE[0].RAM8.WEBUF[1].X ;
 wire \SLICE[0].RAM8.WEBUF[2].A ;
 wire \SLICE[0].RAM8.WEBUF[2].X ;
 wire \SLICE[0].RAM8.WEBUF[3].A ;
 wire \SLICE[0].RAM8.WEBUF[3].X ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[0].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[1].RAM8.CLKBUF.X ;
 wire \SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[1].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[1].RAM8.DEC0.EN ;
 wire \SLICE[1].RAM8.DEC0.EN_buf ;
 wire \SLICE[1].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[1].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[1].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[1].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[1].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[1].RAM8.DEC1.EN ;
 wire \SLICE[1].RAM8.DEC1.EN_buf ;
 wire \SLICE[1].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[1].RAM8.WEBUF[0].X ;
 wire \SLICE[1].RAM8.WEBUF[1].X ;
 wire \SLICE[1].RAM8.WEBUF[2].X ;
 wire \SLICE[1].RAM8.WEBUF[3].X ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[1].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[2].RAM8.CLKBUF.X ;
 wire \SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[2].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[2].RAM8.DEC0.EN ;
 wire \SLICE[2].RAM8.DEC0.EN_buf ;
 wire \SLICE[2].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[2].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[2].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[2].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[2].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[2].RAM8.DEC1.EN ;
 wire \SLICE[2].RAM8.DEC1.EN_buf ;
 wire \SLICE[2].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[2].RAM8.WEBUF[0].X ;
 wire \SLICE[2].RAM8.WEBUF[1].X ;
 wire \SLICE[2].RAM8.WEBUF[2].X ;
 wire \SLICE[2].RAM8.WEBUF[3].X ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[2].RAM8.WORD[7].W.SEL1 ;
 wire \SLICE[3].RAM8.CLKBUF.X ;
 wire \SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC0.A_buf_N[0] ;
 wire \SLICE[3].RAM8.DEC0.A_buf_N[1] ;
 wire \SLICE[3].RAM8.DEC0.EN ;
 wire \SLICE[3].RAM8.DEC0.EN_buf ;
 wire \SLICE[3].RAM8.DEC0.EN_buf_N ;
 wire \SLICE[3].RAM8.DEC1.A_buf[0] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[1] ;
 wire \SLICE[3].RAM8.DEC1.A_buf[2] ;
 wire \SLICE[3].RAM8.DEC1.A_buf_N[0] ;
 wire \SLICE[3].RAM8.DEC1.A_buf_N[1] ;
 wire \SLICE[3].RAM8.DEC1.EN ;
 wire \SLICE[3].RAM8.DEC1.EN_buf ;
 wire \SLICE[3].RAM8.DEC1.EN_buf_N ;
 wire \SLICE[3].RAM8.WEBUF[0].X ;
 wire \SLICE[3].RAM8.WEBUF[1].X ;
 wire \SLICE[3].RAM8.WEBUF[2].X ;
 wire \SLICE[3].RAM8.WEBUF[3].X ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[0].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[1].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[2].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[3].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[4].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[5].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[6].W.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ;
 wire \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \SLICE[3].RAM8.WORD[7].W.SEL1 ;
 wire zero_;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[0].__cell__  (.I(A0[0]),
    .Z(\A0BUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[1].__cell__  (.I(A0[1]),
    .Z(\A0BUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[2].__cell__  (.I(A0[2]),
    .Z(\A0BUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[3].__cell__  (.I(A0[3]),
    .Z(\A0BUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A0BUF[4].__cell__  (.I(A0[4]),
    .Z(\A0BUF[4].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[0].__cell__  (.I(A1[0]),
    .Z(\A1BUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[1].__cell__  (.I(A1[1]),
    .Z(\A1BUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[2].__cell__  (.I(A1[2]),
    .Z(\A1BUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[3].__cell__  (.I(A1[3]),
    .Z(\A1BUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \A1BUF[4].__cell__  (.I(A1[4]),
    .Z(\A1BUF[4].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[0].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[0].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[0].__cell__  (.EN(\BYTE[0].FLOATBUF0[0].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[1].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[1].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[1].__cell__  (.EN(\BYTE[0].FLOATBUF0[1].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[2].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[2].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[2].__cell__  (.EN(\BYTE[0].FLOATBUF0[2].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[3].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[3].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[3].__cell__  (.EN(\BYTE[0].FLOATBUF0[3].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[4].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[4].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[4].__cell__  (.EN(\BYTE[0].FLOATBUF0[4].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[5].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[5].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[5].__cell__  (.EN(\BYTE[0].FLOATBUF0[5].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[6].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[6].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[6].__cell__  (.EN(\BYTE[0].FLOATBUF0[6].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF0[7].TE_BINV  (.I(\BYTE[0].FLOATBUF0[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF0[7].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF0[7].__cell__  (.EN(\BYTE[0].FLOATBUF0[7].TE_BN ),
    .I(\BYTE[0].FLOATBUF0[0].A ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[0].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[0].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[0].__cell__  (.EN(\BYTE[0].FLOATBUF1[0].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[1].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[1].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[1].__cell__  (.EN(\BYTE[0].FLOATBUF1[1].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[2].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[2].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[2].__cell__  (.EN(\BYTE[0].FLOATBUF1[2].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[3].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[3].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[3].__cell__  (.EN(\BYTE[0].FLOATBUF1[3].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[4].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[4].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[4].__cell__  (.EN(\BYTE[0].FLOATBUF1[4].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[5].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[5].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[5].__cell__  (.EN(\BYTE[0].FLOATBUF1[5].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[6].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[6].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[6].__cell__  (.EN(\BYTE[0].FLOATBUF1[6].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[0].FLOATBUF1[7].TE_BINV  (.I(\BYTE[0].FLOATBUF1[0].TE_B ),
    .ZN(\BYTE[0].FLOATBUF1[7].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[0].FLOATBUF1[7].__cell__  (.EN(\BYTE[0].FLOATBUF1[7].TE_BN ),
    .I(\BYTE[0].FLOATBUF1[0].A ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[10].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[10].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[10].__cell__  (.EN(\BYTE[1].FLOATBUF0[10].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[11].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[11].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[11].__cell__  (.EN(\BYTE[1].FLOATBUF0[11].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[12].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[12].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[12].__cell__  (.EN(\BYTE[1].FLOATBUF0[12].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[13].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[13].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[13].__cell__  (.EN(\BYTE[1].FLOATBUF0[13].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[14].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[14].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[14].__cell__  (.EN(\BYTE[1].FLOATBUF0[14].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[15].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[15].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[15].__cell__  (.EN(\BYTE[1].FLOATBUF0[15].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[8].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[8].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[8].__cell__  (.EN(\BYTE[1].FLOATBUF0[8].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF0[9].TE_BINV  (.I(\BYTE[1].FLOATBUF0[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF0[9].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF0[9].__cell__  (.EN(\BYTE[1].FLOATBUF0[9].TE_BN ),
    .I(\BYTE[1].FLOATBUF0[10].A ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[10].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[10].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[10].__cell__  (.EN(\BYTE[1].FLOATBUF1[10].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[11].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[11].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[11].__cell__  (.EN(\BYTE[1].FLOATBUF1[11].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[12].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[12].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[12].__cell__  (.EN(\BYTE[1].FLOATBUF1[12].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[13].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[13].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[13].__cell__  (.EN(\BYTE[1].FLOATBUF1[13].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[14].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[14].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[14].__cell__  (.EN(\BYTE[1].FLOATBUF1[14].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[15].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[15].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[15].__cell__  (.EN(\BYTE[1].FLOATBUF1[15].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[8].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[8].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[8].__cell__  (.EN(\BYTE[1].FLOATBUF1[8].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[1].FLOATBUF1[9].TE_BINV  (.I(\BYTE[1].FLOATBUF1[10].TE_B ),
    .ZN(\BYTE[1].FLOATBUF1[9].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[1].FLOATBUF1[9].__cell__  (.EN(\BYTE[1].FLOATBUF1[9].TE_BN ),
    .I(\BYTE[1].FLOATBUF1[10].A ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[16].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[16].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[16].__cell__  (.EN(\BYTE[2].FLOATBUF0[16].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[17].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[17].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[17].__cell__  (.EN(\BYTE[2].FLOATBUF0[17].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[18].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[18].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[18].__cell__  (.EN(\BYTE[2].FLOATBUF0[18].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[19].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[19].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[19].__cell__  (.EN(\BYTE[2].FLOATBUF0[19].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[20].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[20].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[20].__cell__  (.EN(\BYTE[2].FLOATBUF0[20].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[21].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[21].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[21].__cell__  (.EN(\BYTE[2].FLOATBUF0[21].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[22].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[22].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[22].__cell__  (.EN(\BYTE[2].FLOATBUF0[22].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF0[23].TE_BINV  (.I(\BYTE[2].FLOATBUF0[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF0[23].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF0[23].__cell__  (.EN(\BYTE[2].FLOATBUF0[23].TE_BN ),
    .I(\BYTE[2].FLOATBUF0[16].A ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[16].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[16].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[16].__cell__  (.EN(\BYTE[2].FLOATBUF1[16].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[17].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[17].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[17].__cell__  (.EN(\BYTE[2].FLOATBUF1[17].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[18].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[18].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[18].__cell__  (.EN(\BYTE[2].FLOATBUF1[18].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[19].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[19].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[19].__cell__  (.EN(\BYTE[2].FLOATBUF1[19].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[20].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[20].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[20].__cell__  (.EN(\BYTE[2].FLOATBUF1[20].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[21].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[21].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[21].__cell__  (.EN(\BYTE[2].FLOATBUF1[21].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[22].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[22].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[22].__cell__  (.EN(\BYTE[2].FLOATBUF1[22].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[2].FLOATBUF1[23].TE_BINV  (.I(\BYTE[2].FLOATBUF1[16].TE_B ),
    .ZN(\BYTE[2].FLOATBUF1[23].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[2].FLOATBUF1[23].__cell__  (.EN(\BYTE[2].FLOATBUF1[23].TE_BN ),
    .I(\BYTE[2].FLOATBUF1[16].A ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[24].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[24].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[24].__cell__  (.EN(\BYTE[3].FLOATBUF0[24].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[25].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[25].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[25].__cell__  (.EN(\BYTE[3].FLOATBUF0[25].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[26].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[26].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[26].__cell__  (.EN(\BYTE[3].FLOATBUF0[26].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[27].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[27].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[27].__cell__  (.EN(\BYTE[3].FLOATBUF0[27].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[28].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[28].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[28].__cell__  (.EN(\BYTE[3].FLOATBUF0[28].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[29].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[29].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[29].__cell__  (.EN(\BYTE[3].FLOATBUF0[29].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[30].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[30].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[30].__cell__  (.EN(\BYTE[3].FLOATBUF0[30].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF0[31].TE_BINV  (.I(\BYTE[3].FLOATBUF0[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF0[31].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF0[31].__cell__  (.EN(\BYTE[3].FLOATBUF0[31].TE_BN ),
    .I(\BYTE[3].FLOATBUF0[24].A ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[24].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[24].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[24].__cell__  (.EN(\BYTE[3].FLOATBUF1[24].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[25].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[25].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[25].__cell__  (.EN(\BYTE[3].FLOATBUF1[25].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[26].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[26].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[26].__cell__  (.EN(\BYTE[3].FLOATBUF1[26].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[27].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[27].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[27].__cell__  (.EN(\BYTE[3].FLOATBUF1[27].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[28].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[28].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[28].__cell__  (.EN(\BYTE[3].FLOATBUF1[28].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[29].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[29].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[29].__cell__  (.EN(\BYTE[3].FLOATBUF1[29].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[30].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[30].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[30].__cell__  (.EN(\BYTE[3].FLOATBUF1[30].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \BYTE[3].FLOATBUF1[31].TE_BINV  (.I(\BYTE[3].FLOATBUF1[24].TE_B ),
    .ZN(\BYTE[3].FLOATBUF1[31].TE_BN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \BYTE[3].FLOATBUF1[31].__cell__  (.EN(\BYTE[3].FLOATBUF1[31].TE_BN ),
    .I(\BYTE[3].FLOATBUF1[24].A ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \CLKBUF.__cell__  (.I(CLK),
    .Z(\CLKBUF.X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 \DEC0.AND0  (.A1(\A0BUF[3].X ),
    .A2(\A0BUF[4].X ),
    .A3(\DEC0.EN_N ),
    .ZN(\SLICE[0].RAM8.DEC0.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND1  (.A1(\DEC0.A_N[1] ),
    .A2(\A0BUF[3].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[1].RAM8.DEC0.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND2  (.A1(\DEC0.A_N[0] ),
    .A2(\A0BUF[4].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[2].RAM8.DEC0.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC0.AND3  (.A1(\A0BUF[4].X ),
    .A2(\A0BUF[3].X ),
    .A3(\DEC0.EN ),
    .Z(\SLICE[3].RAM8.DEC0.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV1  (.I(\A0BUF[3].X ),
    .ZN(\DEC0.A_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV2  (.I(\A0BUF[4].X ),
    .ZN(\DEC0.A_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC0.INV3  (.I(\DEC0.EN ),
    .ZN(\DEC0.EN_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 \DEC1.AND0  (.A1(\A1BUF[3].X ),
    .A2(\A1BUF[4].X ),
    .A3(\DEC1.EN_N ),
    .ZN(\SLICE[0].RAM8.DEC1.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND1  (.A1(\DEC1.A_N[1] ),
    .A2(\A1BUF[3].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[1].RAM8.DEC1.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND2  (.A1(\DEC1.A_N[0] ),
    .A2(\A1BUF[4].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[2].RAM8.DEC1.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 \DEC1.AND3  (.A1(\A1BUF[4].X ),
    .A2(\A1BUF[3].X ),
    .A3(\DEC1.EN ),
    .Z(\SLICE[3].RAM8.DEC1.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV1  (.I(\A1BUF[3].X ),
    .ZN(\DEC1.A_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV2  (.I(\A1BUF[4].X ),
    .ZN(\DEC1.A_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \DEC1.INV3  (.I(\DEC1.EN ),
    .ZN(\DEC1.EN_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[0].__cell__  (.I(Di0[0]),
    .Z(\DIBUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[10].__cell__  (.I(Di0[10]),
    .Z(\DIBUF[10].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[11].__cell__  (.I(Di0[11]),
    .Z(\DIBUF[11].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[12].__cell__  (.I(Di0[12]),
    .Z(\DIBUF[12].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[13].__cell__  (.I(Di0[13]),
    .Z(\DIBUF[13].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[14].__cell__  (.I(Di0[14]),
    .Z(\DIBUF[14].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[15].__cell__  (.I(Di0[15]),
    .Z(\DIBUF[15].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[16].__cell__  (.I(Di0[16]),
    .Z(\DIBUF[16].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[17].__cell__  (.I(Di0[17]),
    .Z(\DIBUF[17].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[18].__cell__  (.I(Di0[18]),
    .Z(\DIBUF[18].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[19].__cell__  (.I(Di0[19]),
    .Z(\DIBUF[19].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[1].__cell__  (.I(Di0[1]),
    .Z(\DIBUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[20].__cell__  (.I(Di0[20]),
    .Z(\DIBUF[20].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[21].__cell__  (.I(Di0[21]),
    .Z(\DIBUF[21].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[22].__cell__  (.I(Di0[22]),
    .Z(\DIBUF[22].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[23].__cell__  (.I(Di0[23]),
    .Z(\DIBUF[23].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[24].__cell__  (.I(Di0[24]),
    .Z(\DIBUF[24].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[25].__cell__  (.I(Di0[25]),
    .Z(\DIBUF[25].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[26].__cell__  (.I(Di0[26]),
    .Z(\DIBUF[26].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[27].__cell__  (.I(Di0[27]),
    .Z(\DIBUF[27].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[28].__cell__  (.I(Di0[28]),
    .Z(\DIBUF[28].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[29].__cell__  (.I(Di0[29]),
    .Z(\DIBUF[29].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[2].__cell__  (.I(Di0[2]),
    .Z(\DIBUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[30].__cell__  (.I(Di0[30]),
    .Z(\DIBUF[30].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[31].__cell__  (.I(Di0[31]),
    .Z(\DIBUF[31].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[3].__cell__  (.I(Di0[3]),
    .Z(\DIBUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[4].__cell__  (.I(Di0[4]),
    .Z(\DIBUF[4].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[5].__cell__  (.I(Di0[5]),
    .Z(\DIBUF[5].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[6].__cell__  (.I(Di0[6]),
    .Z(\DIBUF[6].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[7].__cell__  (.I(Di0[7]),
    .Z(\DIBUF[7].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[8].__cell__  (.I(Di0[8]),
    .Z(\DIBUF[8].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \DIBUF[9].__cell__  (.I(Di0[9]),
    .Z(\DIBUF[9].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[0]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[1]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[2]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Do_CLKBUF[3]  (.I(\Do0_REG.CLK_buf ),
    .Z(\Do0_REG.CLKBUF[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.I(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.I(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.I(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.I(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.I(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.I(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.I(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.I(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.D(\BYTE[0].FLOATBUF0[0].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.D(\BYTE[0].FLOATBUF0[1].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.D(\BYTE[0].FLOATBUF0[2].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.D(\BYTE[0].FLOATBUF0[3].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.D(\BYTE[0].FLOATBUF0[4].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.D(\BYTE[0].FLOATBUF0[5].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.D(\BYTE[0].FLOATBUF0[6].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.D(\BYTE[0].FLOATBUF0[7].Z ),
    .CLK(\Do0_REG.CLKBUF[0] ),
    .Q(Do0[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.I(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.I(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.I(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.I(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.I(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.I(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.I(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.I(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.D(\BYTE[1].FLOATBUF0[8].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.D(\BYTE[1].FLOATBUF0[9].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.D(\BYTE[1].FLOATBUF0[10].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.D(\BYTE[1].FLOATBUF0[11].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.D(\BYTE[1].FLOATBUF0[12].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.D(\BYTE[1].FLOATBUF0[13].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.D(\BYTE[1].FLOATBUF0[14].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.D(\BYTE[1].FLOATBUF0[15].Z ),
    .CLK(\Do0_REG.CLKBUF[1] ),
    .Q(Do0[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.I(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.I(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.I(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.I(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.I(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.I(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.I(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.I(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.D(\BYTE[2].FLOATBUF0[16].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.D(\BYTE[2].FLOATBUF0[17].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.D(\BYTE[2].FLOATBUF0[18].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.D(\BYTE[2].FLOATBUF0[19].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.D(\BYTE[2].FLOATBUF0[20].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[20]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.D(\BYTE[2].FLOATBUF0[21].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[21]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.D(\BYTE[2].FLOATBUF0[22].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[22]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.D(\BYTE[2].FLOATBUF0[23].Z ),
    .CLK(\Do0_REG.CLKBUF[2] ),
    .Q(Do0[23]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.I(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.I(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.I(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.I(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.I(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.I(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.I(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.I(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.D(\BYTE[3].FLOATBUF0[24].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[24]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.D(\BYTE[3].FLOATBUF0[25].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[25]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.D(\BYTE[3].FLOATBUF0[26].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[26]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.D(\BYTE[3].FLOATBUF0[27].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[27]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.D(\BYTE[3].FLOATBUF0[28].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[28]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.D(\BYTE[3].FLOATBUF0[29].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[29]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.D(\BYTE[3].FLOATBUF0[30].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[30]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.D(\BYTE[3].FLOATBUF0[31].Z ),
    .CLK(\Do0_REG.CLKBUF[3] ),
    .Q(Do0[31]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do0_REG.Root_CLKBUF  (.I(\CLKBUF.X ),
    .Z(\Do0_REG.CLK_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[0]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[1]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[2]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Do_CLKBUF[3]  (.I(\Do1_REG.CLK_buf ),
    .Z(\Do1_REG.CLKBUF[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[0]  (.I(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[1]  (.I(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[2]  (.I(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[3]  (.I(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[4]  (.I(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[5]  (.I(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[6]  (.I(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[0].DIODE[7]  (.I(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[0]  (.D(\BYTE[0].FLOATBUF1[0].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[1]  (.D(\BYTE[0].FLOATBUF1[1].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[2]  (.D(\BYTE[0].FLOATBUF1[2].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[3]  (.D(\BYTE[0].FLOATBUF1[3].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[4]  (.D(\BYTE[0].FLOATBUF1[4].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[5]  (.D(\BYTE[0].FLOATBUF1[5].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[6]  (.D(\BYTE[0].FLOATBUF1[6].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[0].Do_FF[7]  (.D(\BYTE[0].FLOATBUF1[7].Z ),
    .CLK(\Do1_REG.CLKBUF[0] ),
    .Q(Do1[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[0]  (.I(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[1]  (.I(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[2]  (.I(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[3]  (.I(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[4]  (.I(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[5]  (.I(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[6]  (.I(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[1].DIODE[7]  (.I(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[0]  (.D(\BYTE[1].FLOATBUF1[8].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[1]  (.D(\BYTE[1].FLOATBUF1[9].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[2]  (.D(\BYTE[1].FLOATBUF1[10].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[3]  (.D(\BYTE[1].FLOATBUF1[11].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[4]  (.D(\BYTE[1].FLOATBUF1[12].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[5]  (.D(\BYTE[1].FLOATBUF1[13].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[6]  (.D(\BYTE[1].FLOATBUF1[14].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[1].Do_FF[7]  (.D(\BYTE[1].FLOATBUF1[15].Z ),
    .CLK(\Do1_REG.CLKBUF[1] ),
    .Q(Do1[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[0]  (.I(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[1]  (.I(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[2]  (.I(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[3]  (.I(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[4]  (.I(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[5]  (.I(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[6]  (.I(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[2].DIODE[7]  (.I(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[0]  (.D(\BYTE[2].FLOATBUF1[16].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[1]  (.D(\BYTE[2].FLOATBUF1[17].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[2]  (.D(\BYTE[2].FLOATBUF1[18].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[3]  (.D(\BYTE[2].FLOATBUF1[19].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[4]  (.D(\BYTE[2].FLOATBUF1[20].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[20]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[5]  (.D(\BYTE[2].FLOATBUF1[21].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[21]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[6]  (.D(\BYTE[2].FLOATBUF1[22].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[22]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[2].Do_FF[7]  (.D(\BYTE[2].FLOATBUF1[23].Z ),
    .CLK(\Do1_REG.CLKBUF[2] ),
    .Q(Do1[23]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[0]  (.I(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[1]  (.I(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[2]  (.I(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[3]  (.I(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[4]  (.I(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[5]  (.I(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[6]  (.I(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \Do1_REG.OUTREG_BYTE[3].DIODE[7]  (.I(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[0]  (.D(\BYTE[3].FLOATBUF1[24].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[24]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[1]  (.D(\BYTE[3].FLOATBUF1[25].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[25]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[2]  (.D(\BYTE[3].FLOATBUF1[26].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[26]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[3]  (.D(\BYTE[3].FLOATBUF1[27].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[27]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[4]  (.D(\BYTE[3].FLOATBUF1[28].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[28]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[5]  (.D(\BYTE[3].FLOATBUF1[29].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[29]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[6]  (.D(\BYTE[3].FLOATBUF1[30].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[30]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \Do1_REG.OUTREG_BYTE[3].Do_FF[7]  (.D(\BYTE[3].FLOATBUF1[31].Z ),
    .CLK(\Do1_REG.CLKBUF[3] ),
    .Q(Do1[31]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \Do1_REG.Root_CLKBUF  (.I(\CLKBUF.X ),
    .Z(\Do1_REG.CLK_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \EN0BUF.__cell__  (.I(EN0),
    .Z(\DEC0.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \EN1BUF.__cell__  (.I(EN1),
    .Z(\DEC1.EN ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[0].__cell__  (.I(EN0),
    .Z(\BYTE[0].FLOATBUF0[0].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[1].__cell__  (.I(EN0),
    .Z(\BYTE[1].FLOATBUF0[10].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[2].__cell__  (.I(EN0),
    .Z(\BYTE[2].FLOATBUF0[16].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF0[3].__cell__  (.I(EN0),
    .Z(\BYTE[3].FLOATBUF0[24].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[0].__cell__  (.I(EN1),
    .Z(\BYTE[0].FLOATBUF1[0].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[1].__cell__  (.I(EN1),
    .Z(\BYTE[1].FLOATBUF1[10].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[2].__cell__  (.I(EN1),
    .Z(\BYTE[2].FLOATBUF1[16].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \FBUFENBUF1[3].__cell__  (.I(EN1),
    .Z(\BYTE[3].FLOATBUF1[24].TE_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[0].RAM8.CLKBUF.X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[0].RAM8.DEC0.AND0  (.A1(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND4  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND5  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND6  (.A1(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC0.AND7  (.A1(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC0.ENBUF  (.I(\SLICE[0].RAM8.DEC0.EN ),
    .Z(\SLICE[0].RAM8.DEC0.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV1  (.I(\SLICE[0].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV2  (.I(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV3  (.I(\SLICE[0].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC0.INV4  (.I(\SLICE[0].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[0].RAM8.DEC0.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[0].RAM8.DEC1.AND0  (.A1(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[1].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[2].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[3].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND4  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[4].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND5  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[5].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND6  (.A1(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[6].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[0].RAM8.DEC1.AND7  (.A1(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[0].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[0].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[0].RAM8.WORD[7].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.DEC1.ENBUF  (.I(\SLICE[0].RAM8.DEC1.EN ),
    .Z(\SLICE[0].RAM8.DEC1.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV1  (.I(\SLICE[0].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV2  (.I(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV3  (.I(\SLICE[0].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[0].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.DEC1.INV4  (.I(\SLICE[0].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[0].RAM8.DEC1.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[0].RAM8.WEBUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[0].RAM8.WEBUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[0].RAM8.WEBUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[0].RAM8.WEBUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[0].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[1].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[2].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[0].RAM8.WEBUF[3].X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[0].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[0].RAM8.CLKBUF.X ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[0].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[0].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[1].RAM8.CLKBUF.X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[1].RAM8.DEC0.AND0  (.A1(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND4  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND5  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND6  (.A1(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC0.AND7  (.A1(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC0.ENBUF  (.I(\SLICE[1].RAM8.DEC0.EN ),
    .Z(\SLICE[1].RAM8.DEC0.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV1  (.I(\SLICE[1].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV2  (.I(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV3  (.I(\SLICE[1].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC0.INV4  (.I(\SLICE[1].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[1].RAM8.DEC0.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[1].RAM8.DEC1.AND0  (.A1(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[1].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[2].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[3].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND4  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[4].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND5  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[5].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND6  (.A1(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[6].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[1].RAM8.DEC1.AND7  (.A1(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[1].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[1].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[1].RAM8.WORD[7].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.DEC1.ENBUF  (.I(\SLICE[1].RAM8.DEC1.EN ),
    .Z(\SLICE[1].RAM8.DEC1.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV1  (.I(\SLICE[1].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV2  (.I(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV3  (.I(\SLICE[1].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[1].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.DEC1.INV4  (.I(\SLICE[1].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[1].RAM8.DEC1.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[1].RAM8.WEBUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[1].RAM8.WEBUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[1].RAM8.WEBUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[1].RAM8.WEBUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[0].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[1].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[2].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[1].RAM8.WEBUF[3].X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[1].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[1].RAM8.CLKBUF.X ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[1].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[1].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[2].RAM8.CLKBUF.X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[2].RAM8.DEC0.AND0  (.A1(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND4  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND5  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND6  (.A1(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC0.AND7  (.A1(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC0.ENBUF  (.I(\SLICE[2].RAM8.DEC0.EN ),
    .Z(\SLICE[2].RAM8.DEC0.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV1  (.I(\SLICE[2].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV2  (.I(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV3  (.I(\SLICE[2].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC0.INV4  (.I(\SLICE[2].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[2].RAM8.DEC0.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[2].RAM8.DEC1.AND0  (.A1(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[1].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[2].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[3].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND4  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[4].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND5  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[5].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND6  (.A1(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[6].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[2].RAM8.DEC1.AND7  (.A1(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[2].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[2].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[2].RAM8.WORD[7].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.DEC1.ENBUF  (.I(\SLICE[2].RAM8.DEC1.EN ),
    .Z(\SLICE[2].RAM8.DEC1.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV1  (.I(\SLICE[2].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV2  (.I(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV3  (.I(\SLICE[2].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[2].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.DEC1.INV4  (.I(\SLICE[2].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[2].RAM8.DEC1.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[2].RAM8.WEBUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[2].RAM8.WEBUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[2].RAM8.WEBUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[2].RAM8.WEBUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[0].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[1].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[2].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[2].RAM8.WEBUF[3].X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[2].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[2].RAM8.CLKBUF.X ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[2].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[2].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.CLKBUF.__cell__  (.I(\CLKBUF.X ),
    .Z(\SLICE[3].RAM8.CLKBUF.X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[0]  (.I(\A0BUF[0].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[1]  (.I(\A0BUF[1].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ABUF[2]  (.I(\A0BUF[2].X ),
    .Z(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[3].RAM8.DEC0.AND0  (.A1(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf_N ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND1  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND2  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND3  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND4  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND5  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND6  (.A1(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC0.AND7  (.A1(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC0.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC0.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC0.ENBUF  (.I(\SLICE[3].RAM8.DEC0.EN ),
    .Z(\SLICE[3].RAM8.DEC0.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV1  (.I(\SLICE[3].RAM8.DEC0.A_buf[0] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV2  (.I(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV3  (.I(\SLICE[3].RAM8.DEC0.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC0.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC0.INV4  (.I(\SLICE[3].RAM8.DEC0.EN_buf ),
    .ZN(\SLICE[3].RAM8.DEC0.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[0]  (.I(\A1BUF[0].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[1]  (.I(\A1BUF[1].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ABUF[2]  (.I(\A1BUF[2].X ),
    .Z(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \SLICE[3].RAM8.DEC1.AND0  (.A1(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf_N ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND1  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[1].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND2  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[2].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND3  (.A1(zero_),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[3].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND4  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[4].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND5  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[5].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND6  (.A1(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[6].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 \SLICE[3].RAM8.DEC1.AND7  (.A1(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .A2(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .A3(\SLICE[3].RAM8.DEC1.A_buf[2] ),
    .A4(\SLICE[3].RAM8.DEC1.EN_buf ),
    .Z(\SLICE[3].RAM8.WORD[7].W.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.DEC1.ENBUF  (.I(\SLICE[3].RAM8.DEC1.EN ),
    .Z(\SLICE[3].RAM8.DEC1.EN_buf ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV1  (.I(\SLICE[3].RAM8.DEC1.A_buf[0] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV2  (.I(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV3  (.I(\SLICE[3].RAM8.DEC1.A_buf[1] ),
    .ZN(\SLICE[3].RAM8.DEC1.A_buf_N[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.DEC1.INV4  (.I(\SLICE[3].RAM8.DEC1.EN_buf ),
    .ZN(\SLICE[3].RAM8.DEC1.EN_buf_N ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[0].__cell__  (.I(\SLICE[0].RAM8.WEBUF[0].A ),
    .Z(\SLICE[3].RAM8.WEBUF[0].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[1].__cell__  (.I(\SLICE[0].RAM8.WEBUF[1].A ),
    .Z(\SLICE[3].RAM8.WEBUF[1].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[2].__cell__  (.I(\SLICE[0].RAM8.WEBUF[2].A ),
    .Z(\SLICE[3].RAM8.WEBUF[2].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WEBUF[3].__cell__  (.I(\SLICE[0].RAM8.WEBUF[3].A ),
    .Z(\SLICE[3].RAM8.WEBUF[3].X ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[0].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[0].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[0].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[1].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[1].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[1].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[2].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[2].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[2].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[3].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[3].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[3].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[4].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[4].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[4].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[5].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[5].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[5].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[6].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[6].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[6].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF0[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .Z(\BYTE[0].FLOATBUF1[0].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[0].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF0[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .Z(\BYTE[0].FLOATBUF1[1].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[1].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF0[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .Z(\BYTE[0].FLOATBUF1[2].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[2].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF0[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .Z(\BYTE[0].FLOATBUF1[3].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[3].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF0[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .Z(\BYTE[0].FLOATBUF1[4].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[4].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF0[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .Z(\BYTE[0].FLOATBUF1[5].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[5].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF0[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .Z(\BYTE[0].FLOATBUF1[6].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[6].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF0[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .Z(\BYTE[0].FLOATBUF1[7].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[7].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[0].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF0[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .Z(\BYTE[1].FLOATBUF1[8].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[8].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF0[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .Z(\BYTE[1].FLOATBUF1[9].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[9].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF0[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .Z(\BYTE[1].FLOATBUF1[10].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[10].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF0[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .Z(\BYTE[1].FLOATBUF1[11].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[11].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF0[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .Z(\BYTE[1].FLOATBUF1[12].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[12].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF0[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .Z(\BYTE[1].FLOATBUF1[13].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[13].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF0[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .Z(\BYTE[1].FLOATBUF1[14].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[14].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF0[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .Z(\BYTE[1].FLOATBUF1[15].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[15].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[1].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF0[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .Z(\BYTE[2].FLOATBUF1[16].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[16].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF0[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .Z(\BYTE[2].FLOATBUF1[17].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[17].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF0[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .Z(\BYTE[2].FLOATBUF1[18].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[18].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF0[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .Z(\BYTE[2].FLOATBUF1[19].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[19].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF0[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .Z(\BYTE[2].FLOATBUF1[20].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[20].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF0[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .Z(\BYTE[2].FLOATBUF1[21].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[21].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF0[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .Z(\BYTE[2].FLOATBUF1[22].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[22].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF0[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .Z(\BYTE[2].FLOATBUF1[23].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[23].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[2].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF0[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .Z(\BYTE[3].FLOATBUF1[24].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\DIBUF[24].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF0[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .Z(\BYTE[3].FLOATBUF1[25].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\DIBUF[25].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF0[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .Z(\BYTE[3].FLOATBUF1[26].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\DIBUF[26].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF0[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .Z(\BYTE[3].FLOATBUF1[27].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\DIBUF[27].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF0[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .Z(\BYTE[3].FLOATBUF1[28].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\DIBUF[28].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF0[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .Z(\BYTE[3].FLOATBUF1[29].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\DIBUF[29].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF0[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .Z(\BYTE[3].FLOATBUF1[30].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\DIBUF[30].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF0[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__bufz_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF1  (.EN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .I(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .Z(\BYTE[3].FLOATBUF1[31].Z ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\DIBUF[31].X ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A1(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .A2(\SLICE[3].RAM8.WEBUF[3].X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1INV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL1_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__icgtp_1 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .E(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .TE(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .Q(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.I(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .ZN(\SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \SLICE[3].RAM8.WORD[7].W.CLKBUF  (.I(\SLICE[3].RAM8.CLKBUF.X ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.I(\SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \SLICE[3].RAM8.WORD[7].W.SEL1BUF  (.I(\SLICE[3].RAM8.WORD[7].W.SEL1 ),
    .Z(\SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[0].__cell__  (.ZN(\BYTE[0].FLOATBUF0[0].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[1].__cell__  (.ZN(\BYTE[1].FLOATBUF0[10].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[2].__cell__  (.ZN(\BYTE[2].FLOATBUF0[16].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE0[3].__cell__  (.ZN(\BYTE[3].FLOATBUF0[24].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[0].__cell__  (.ZN(\BYTE[0].FLOATBUF1[0].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[1].__cell__  (.ZN(\BYTE[1].FLOATBUF1[10].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[2].__cell__  (.ZN(\BYTE[2].FLOATBUF1[16].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel \TIE1[3].__cell__  (.ZN(\BYTE[3].FLOATBUF1[24].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[0].__cell__  (.I(WE0[0]),
    .Z(\SLICE[0].RAM8.WEBUF[0].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[1].__cell__  (.I(WE0[1]),
    .Z(\SLICE[0].RAM8.WEBUF[1].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[2].__cell__  (.I(WE0[2]),
    .Z(\SLICE[0].RAM8.WEBUF[2].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \WEBUF[3].__cell__  (.I(WE0[3]),
    .Z(\SLICE[0].RAM8.WEBUF[3].A ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__tiel TIE_ZERO_zero_ (.ZN(zero_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_0_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_1_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_2_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_3_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_4_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_13_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_15_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_5_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_7_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_8_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_2_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_3_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_4_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_5_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_6_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_6_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_7_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_7_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_8_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_6_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_7_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_8_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_1_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_2_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_4_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_13_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_13_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_14_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_15_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_15_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_16_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_13_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_14_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_15_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_16_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_9_60 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_10_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_12_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_14_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_15_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_16_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_21_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_23_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_18_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_18_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_19_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_20_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_20_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_21_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_21_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_22_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_22_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_23_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_23_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_24_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_24_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_22_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_23_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_24_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_17_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_18_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_20_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_22_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_24_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_29_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_31_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_26_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_26_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_27_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_28_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_28_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_29_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_29_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_30_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_30_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_31_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_31_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_32_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_32_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_27_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_30_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_31_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_32_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_25_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_26_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_28_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_30_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_32_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_33_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_60 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_61 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_62 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_63 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_64 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_65 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_66 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_67 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_68 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_69 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_34_70 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_0_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_3_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_6_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_11_60 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie tap_19_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_254 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_256 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_258 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_261 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_264 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_270 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_272 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_273 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_275 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_280 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_281 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_283 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_285 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_286 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_287 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_288 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_289 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_291 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_293 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_294 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_295 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_296 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_297 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_298 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_299 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_300 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_301 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_303 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_305 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_306 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_307 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_309 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_310 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_311 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_315 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_316 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_318 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_319 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_320 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_321 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_323 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_324 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_326 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_328 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_330 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_331 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_332 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_333 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_334 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_335 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_336 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_338 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_339 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_340 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_341 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_343 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_344 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_345 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_346 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_347 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_350 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_351 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_353 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_354 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_355 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_356 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_357 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_358 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_359 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_360 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_361 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_363 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_365 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_366 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_367 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_368 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_370 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_371 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_373 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_375 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_376 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_377 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_379 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_380 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_381 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_385 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_386 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_388 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_389 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_390 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_391 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_392 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_393 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_394 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_396 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_397 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_398 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_400 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_402 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_404 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_405 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_406 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_408 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_409 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_410 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_411 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_412 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_413 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_414 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_415 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_416 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_417 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_420 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_421 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_423 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_424 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_425 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_426 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_427 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_428 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_429 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_430 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_431 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_432 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_433 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_434 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_435 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_436 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_438 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_439 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_440 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_441 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_443 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_444 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_445 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_446 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_447 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_448 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_449 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_450 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_451 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_452 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_455 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_456 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_458 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_459 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_460 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_461 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_462 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_463 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_464 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_467 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_470 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_471 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_472 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_473 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_474 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_475 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_476 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_477 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_478 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_479 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_480 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_481 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_482 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_483 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_484 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_486 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_490 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_491 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_493 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_494 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_495 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_499 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_500 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_501 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_502 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_503 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_504 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_505 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_506 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_507 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_508 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_509 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_510 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_511 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_512 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_513 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_514 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_515 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_516 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_517 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_0_518 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_0_519 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_0_520 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_0_521 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_0_522 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_0_523 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_1_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_1_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_1_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_1_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_1_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_1_209 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_2_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_2_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_2_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_2_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_2_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_2_218 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_3_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_3_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_3_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_3_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_3_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_3_216 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_4_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_4_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_4_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_4_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_4_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_4_218 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_5_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_5_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_5_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_5_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_5_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_5_235 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_6_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_6_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_6_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_6_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_6_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_6_225 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_7_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_7_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_7_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_7_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_7_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_7_231 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_8_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_8_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_8_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_8_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_8_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_8_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_9_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_9_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_9_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_9_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_9_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_9_202 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_10_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_10_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_10_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_10_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_10_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_10_220 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_11_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_11_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_11_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_11_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_11_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_11_216 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_12_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_12_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_12_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_12_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_12_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_12_220 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_13_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_13_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_13_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_13_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_13_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_13_231 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_14_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_14_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_14_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_14_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_14_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_14_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_15_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_15_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_15_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_15_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_15_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_15_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_16_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_16_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_16_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_16_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_16_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_16_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_17_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_17_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_17_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_17_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_17_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_17_212 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_18_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_18_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_18_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_18_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_18_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_18_228 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_19_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_19_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_19_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_19_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_19_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_19_225 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_20_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_20_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_20_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_20_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_20_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_20_228 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_21_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_21_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_21_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_21_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_21_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_21_244 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_22_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_22_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_22_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_22_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_22_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_22_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_23_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_23_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_23_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_23_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_23_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_23_253 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_24_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_24_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_24_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_24_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_24_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_24_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_25_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_25_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_25_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_25_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_25_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_25_226 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_26_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_26_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_26_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_26_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_26_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_26_236 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_27_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_27_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_27_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_27_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_27_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_27_235 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_28_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_28_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_28_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_28_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_28_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_28_236 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_29_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_29_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_29_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_29_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_29_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_29_252 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_30_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_30_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_30_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_30_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_30_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_30_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_31_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_31_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_31_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_31_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_31_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_31_253 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_32_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_32_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_32_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_32_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_32_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_32_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_0 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_1 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_3 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_5 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_7 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_9 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_11 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_12 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_15 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_17 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_18 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_19 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_20 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_21 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_28 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_29 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_31 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_36 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_38 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_40 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_42 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_44 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_47 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_50 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_55 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_56 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_58 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_59 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_65 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_66 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_81 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_85 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_88 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_90 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_93 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_94 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_95 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_108 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_110 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_112 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_129 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_135 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_140 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_143 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_145 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_152 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_160 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_188 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_197 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_210 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_215 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_217 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_225 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_229 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_231 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_234 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_235 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_250 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_254 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_256 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_258 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_260 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_261 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_262 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_264 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_270 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_272 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_273 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_275 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_280 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_281 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_283 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_285 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_286 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_287 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_288 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_289 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_291 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_293 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_294 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_295 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_296 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_297 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_298 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_299 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_300 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_301 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_303 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_305 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_306 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_307 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_309 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_310 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_311 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_315 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_316 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_318 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_319 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_320 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_321 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_323 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_324 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_326 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_328 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_330 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_331 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_332 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_333 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_334 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_335 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_336 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_338 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_339 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_340 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_341 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_343 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_344 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_345 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_346 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_347 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_350 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_351 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_353 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_354 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_355 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_356 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_357 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_358 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_359 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_360 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_361 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_363 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_365 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_366 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_367 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_368 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_370 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_371 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_373 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_375 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_376 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_377 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_379 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_380 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_381 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_385 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_386 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_388 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_389 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_390 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_391 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_392 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_393 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_394 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_396 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_397 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_398 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_400 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_402 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_404 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_405 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_406 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_408 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_409 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_410 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_411 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_412 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_413 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_414 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_415 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_416 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_417 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_420 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_421 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_423 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_424 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_425 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_426 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_427 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_428 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_429 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_430 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_431 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_432 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_433 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_434 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_435 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_436 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_438 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_439 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_440 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_441 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_443 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_444 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_445 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_446 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_447 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_448 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_449 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_450 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_451 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_452 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_455 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_456 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_458 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_459 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_460 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_461 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_462 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_463 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_464 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_467 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_470 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_471 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_472 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_473 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_474 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_475 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_476 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_477 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_478 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_479 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_480 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_481 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_482 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_483 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_484 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_486 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_490 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_491 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_493 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_494 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_495 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_499 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_500 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_501 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_502 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_503 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_504 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_505 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_506 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_507 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_508 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_509 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_510 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_511 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_512 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_513 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_514 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_515 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_516 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_517 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_518 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_519 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_520 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_521 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_522 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_523 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_524 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_525 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_526 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_527 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_528 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_529 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_530 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_531 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_532 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_533 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_534 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_535 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_536 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_537 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_538 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_539 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_540 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_541 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_542 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_543 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_544 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_545 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_546 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_547 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_548 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_549 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_550 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_551 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_552 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_553 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_554 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_555 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_556 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_557 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_558 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_559 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_560 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_561 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_562 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_563 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_564 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_565 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_566 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_567 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_568 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_569 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_570 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_571 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_572 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_573 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_574 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_575 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_576 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_577 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_578 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_579 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_580 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_581 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_582 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_583 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_584 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_585 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_586 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_587 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_588 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_589 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_590 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_591 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_592 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_593 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_594 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_595 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_596 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_597 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_598 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_599 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_600 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_601 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_602 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_603 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_604 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_605 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_606 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_607 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_608 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_609 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_610 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_611 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_612 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_613 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_614 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_615 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_616 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_617 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_618 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_619 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_620 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_621 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_622 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_623 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_624 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_625 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_626 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_627 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_628 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_629 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_630 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_631 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_632 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_633 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_634 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_635 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_636 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_637 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_638 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_639 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_640 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_641 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_642 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_643 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_644 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_645 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_646 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_647 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_648 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_649 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_650 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_651 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_652 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_653 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_654 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_655 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_656 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_657 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_658 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_659 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_660 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_661 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_662 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_663 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_664 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_665 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_666 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_667 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_668 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_669 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_670 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_671 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_672 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_673 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_674 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_675 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_676 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_677 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_678 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_679 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_680 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_681 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_682 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_683 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_684 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_685 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_686 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_687 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_688 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_689 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_690 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_691 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_692 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_693 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_694 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_695 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_696 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_697 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_698 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_699 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_700 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_701 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_702 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_703 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_704 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_705 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_706 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_707 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_708 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_709 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_710 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_711 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_712 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_713 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_714 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_715 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_716 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_717 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_718 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_719 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_720 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_721 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_722 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_723 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_724 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_725 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_726 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_727 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_728 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_729 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_730 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_731 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_732 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_733 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_734 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_735 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_736 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_737 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_738 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_739 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_740 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_741 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_742 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_743 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_744 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_745 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_746 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_747 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_748 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_749 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_750 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_751 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_752 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_753 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_754 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_755 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_756 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_757 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_758 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_759 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_760 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_761 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_762 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_763 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_764 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_765 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_766 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_767 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_768 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_769 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_770 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_771 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_772 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_773 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_774 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_775 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_776 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_777 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_778 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_779 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_780 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_781 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_782 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_783 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_784 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_785 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_786 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_787 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_788 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_789 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_790 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_791 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_792 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_793 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_794 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_795 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_796 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 fill_33_797 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 fill_33_798 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 fill_33_799 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 fill_33_800 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 fill_33_801 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie fill_33_802 (.VDD(VDD),
    .VSS(VSS));
endmodule
