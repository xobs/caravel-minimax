// This is the unpowered netlist.
module mimi (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire net359;
 wire net358;
 wire net357;
 wire net356;
 wire net355;
 wire net354;
 wire net353;
 wire net352;
 wire net351;
 wire net350;
 wire net349;
 wire net348;
 wire net347;
 wire net346;
 wire net345;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net385;
 wire net384;
 wire net383;
 wire net382;
 wire net381;
 wire net380;
 wire net379;
 wire net378;
 wire net377;
 wire net376;
 wire net375;
 wire net374;
 wire net373;
 wire net372;
 wire net371;
 wire net370;
 wire net369;
 wire net368;
 wire net367;
 wire net366;
 wire net365;
 wire net364;
 wire \clknet_1_1__leaf_bank1.cen ;
 wire \clknet_1_0__leaf_bank1.cen ;
 wire \clknet_0_bank1.cen ;
 wire \clknet_1_1__leaf_bank2.cen ;
 wire \clknet_1_0__leaf_bank2.cen ;
 wire \clknet_0_bank2.cen ;
 wire \clknet_1_1__leaf_bank3.cen ;
 wire \clknet_1_0__leaf_bank3.cen ;
 wire \clknet_0_bank3.cen ;
 wire \clknet_1_1__leaf_bank4.cen ;
 wire \clknet_1_0__leaf_bank4.cen ;
 wire \clknet_0_bank4.cen ;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_1_1_0_wb_clk_i;
 wire clknet_1_0_0_wb_clk_i;
 wire net363;
 wire net362;
 wire net361;
 wire net169;
 wire \bank1.addr[0] ;
 wire \bank1.addr[1] ;
 wire \bank1.addr[2] ;
 wire \bank1.addr[3] ;
 wire \bank1.addr[4] ;
 wire \bank1.addr[5] ;
 wire \bank1.addr[6] ;
 wire \bank1.addr[7] ;
 wire \bank1.addr[8] ;
 wire \bank1.cen ;
 wire clknet_0_wb_clk_i;
 wire \bank1.rdata[0] ;
 wire \bank1.rdata[10] ;
 wire \bank1.rdata[11] ;
 wire \bank1.rdata[12] ;
 wire \bank1.rdata[13] ;
 wire \bank1.rdata[14] ;
 wire \bank1.rdata[15] ;
 wire \bank1.rdata[16] ;
 wire \bank1.rdata[17] ;
 wire \bank1.rdata[18] ;
 wire \bank1.rdata[19] ;
 wire \bank1.rdata[1] ;
 wire \bank1.rdata[20] ;
 wire \bank1.rdata[21] ;
 wire \bank1.rdata[22] ;
 wire \bank1.rdata[23] ;
 wire \bank1.rdata[24] ;
 wire \bank1.rdata[25] ;
 wire \bank1.rdata[26] ;
 wire \bank1.rdata[27] ;
 wire \bank1.rdata[28] ;
 wire \bank1.rdata[29] ;
 wire \bank1.rdata[2] ;
 wire \bank1.rdata[30] ;
 wire \bank1.rdata[31] ;
 wire \bank1.rdata[3] ;
 wire \bank1.rdata[4] ;
 wire \bank1.rdata[5] ;
 wire \bank1.rdata[6] ;
 wire \bank1.rdata[7] ;
 wire \bank1.rdata[8] ;
 wire \bank1.rdata[9] ;
 wire \bank1.was_en ;
 wire \bank1.wen_mask[0] ;
 wire \bank2.cen ;
 wire \bank2.rdata[0] ;
 wire \bank2.rdata[10] ;
 wire \bank2.rdata[11] ;
 wire \bank2.rdata[12] ;
 wire \bank2.rdata[13] ;
 wire \bank2.rdata[14] ;
 wire \bank2.rdata[15] ;
 wire \bank2.rdata[16] ;
 wire \bank2.rdata[17] ;
 wire \bank2.rdata[18] ;
 wire \bank2.rdata[19] ;
 wire \bank2.rdata[1] ;
 wire \bank2.rdata[20] ;
 wire \bank2.rdata[21] ;
 wire \bank2.rdata[22] ;
 wire \bank2.rdata[23] ;
 wire \bank2.rdata[24] ;
 wire \bank2.rdata[25] ;
 wire \bank2.rdata[26] ;
 wire \bank2.rdata[27] ;
 wire \bank2.rdata[28] ;
 wire \bank2.rdata[29] ;
 wire \bank2.rdata[2] ;
 wire \bank2.rdata[30] ;
 wire \bank2.rdata[31] ;
 wire \bank2.rdata[3] ;
 wire \bank2.rdata[4] ;
 wire \bank2.rdata[5] ;
 wire \bank2.rdata[6] ;
 wire \bank2.rdata[7] ;
 wire \bank2.rdata[8] ;
 wire \bank2.rdata[9] ;
 wire \bank2.was_en ;
 wire \bank3.cen ;
 wire \bank3.rdata[0] ;
 wire \bank3.rdata[10] ;
 wire \bank3.rdata[11] ;
 wire \bank3.rdata[12] ;
 wire \bank3.rdata[13] ;
 wire \bank3.rdata[14] ;
 wire \bank3.rdata[15] ;
 wire \bank3.rdata[16] ;
 wire \bank3.rdata[17] ;
 wire \bank3.rdata[18] ;
 wire \bank3.rdata[19] ;
 wire \bank3.rdata[1] ;
 wire \bank3.rdata[20] ;
 wire \bank3.rdata[21] ;
 wire \bank3.rdata[22] ;
 wire \bank3.rdata[23] ;
 wire \bank3.rdata[24] ;
 wire \bank3.rdata[25] ;
 wire \bank3.rdata[26] ;
 wire \bank3.rdata[27] ;
 wire \bank3.rdata[28] ;
 wire \bank3.rdata[29] ;
 wire \bank3.rdata[2] ;
 wire \bank3.rdata[30] ;
 wire \bank3.rdata[31] ;
 wire \bank3.rdata[3] ;
 wire \bank3.rdata[4] ;
 wire \bank3.rdata[5] ;
 wire \bank3.rdata[6] ;
 wire \bank3.rdata[7] ;
 wire \bank3.rdata[8] ;
 wire \bank3.rdata[9] ;
 wire \bank3.was_en ;
 wire \bank4.cen ;
 wire \bank4.rdata[0] ;
 wire \bank4.rdata[10] ;
 wire \bank4.rdata[11] ;
 wire \bank4.rdata[12] ;
 wire \bank4.rdata[13] ;
 wire \bank4.rdata[14] ;
 wire \bank4.rdata[15] ;
 wire \bank4.rdata[16] ;
 wire \bank4.rdata[17] ;
 wire \bank4.rdata[18] ;
 wire \bank4.rdata[19] ;
 wire \bank4.rdata[1] ;
 wire \bank4.rdata[20] ;
 wire \bank4.rdata[21] ;
 wire \bank4.rdata[22] ;
 wire \bank4.rdata[23] ;
 wire \bank4.rdata[24] ;
 wire \bank4.rdata[25] ;
 wire \bank4.rdata[26] ;
 wire \bank4.rdata[27] ;
 wire \bank4.rdata[28] ;
 wire \bank4.rdata[29] ;
 wire \bank4.rdata[2] ;
 wire \bank4.rdata[30] ;
 wire \bank4.rdata[31] ;
 wire \bank4.rdata[3] ;
 wire \bank4.rdata[4] ;
 wire \bank4.rdata[5] ;
 wire \bank4.rdata[6] ;
 wire \bank4.rdata[7] ;
 wire \bank4.rdata[8] ;
 wire \bank4.rdata[9] ;
 wire \bank4.was_en ;
 wire \inst_lat[0] ;
 wire \inst_lat[10] ;
 wire \inst_lat[11] ;
 wire \inst_lat[12] ;
 wire \inst_lat[13] ;
 wire \inst_lat[14] ;
 wire \inst_lat[15] ;
 wire \inst_lat[1] ;
 wire \inst_lat[2] ;
 wire \inst_lat[3] ;
 wire \inst_lat[4] ;
 wire \inst_lat[5] ;
 wire \inst_lat[6] ;
 wire \inst_lat[7] ;
 wire \inst_lat[8] ;
 wire \inst_lat[9] ;
 wire net170;
 wire net171;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net172;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net173;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net222;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net223;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net213;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net214;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net215;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net216;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net217;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net218;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net219;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net220;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net221;
 wire \minimax.addrD_port[0] ;
 wire \minimax.addrD_port[1] ;
 wire \minimax.addrD_port[2] ;
 wire \minimax.addrD_port[3] ;
 wire \minimax.addrD_port[4] ;
 wire \minimax.addrS_port[0] ;
 wire \minimax.addrS_port[1] ;
 wire \minimax.addrS_port[2] ;
 wire \minimax.addrS_port[3] ;
 wire \minimax.addrS_port[4] ;
 wire \minimax.aluX[0] ;
 wire \minimax.aluX[10] ;
 wire \minimax.aluX[11] ;
 wire \minimax.aluX[12] ;
 wire \minimax.aluX[13] ;
 wire \minimax.aluX[14] ;
 wire \minimax.aluX[15] ;
 wire \minimax.aluX[16] ;
 wire \minimax.aluX[17] ;
 wire \minimax.aluX[18] ;
 wire \minimax.aluX[19] ;
 wire \minimax.aluX[1] ;
 wire \minimax.aluX[20] ;
 wire \minimax.aluX[21] ;
 wire \minimax.aluX[22] ;
 wire \minimax.aluX[23] ;
 wire \minimax.aluX[24] ;
 wire \minimax.aluX[25] ;
 wire \minimax.aluX[26] ;
 wire \minimax.aluX[27] ;
 wire \minimax.aluX[28] ;
 wire \minimax.aluX[29] ;
 wire \minimax.aluX[2] ;
 wire \minimax.aluX[30] ;
 wire \minimax.aluX[31] ;
 wire \minimax.aluX[3] ;
 wire \minimax.aluX[4] ;
 wire \minimax.aluX[5] ;
 wire \minimax.aluX[6] ;
 wire \minimax.aluX[7] ;
 wire \minimax.aluX[8] ;
 wire \minimax.aluX[9] ;
 wire \minimax.bubble1 ;
 wire \minimax.bubble2 ;
 wire \minimax.dly16_lw ;
 wire \minimax.dly16_lwsp ;
 wire \minimax.dly16_slli_setrd ;
 wire \minimax.dly16_slli_setrs ;
 wire \minimax.dra[0] ;
 wire \minimax.dra[1] ;
 wire \minimax.dra[2] ;
 wire \minimax.dra[3] ;
 wire \minimax.dra[4] ;
 wire \minimax.inst[0] ;
 wire \minimax.inst[10] ;
 wire \minimax.inst[11] ;
 wire \minimax.inst[12] ;
 wire \minimax.inst[13] ;
 wire \minimax.inst[14] ;
 wire \minimax.inst[15] ;
 wire \minimax.inst[1] ;
 wire \minimax.inst[2] ;
 wire \minimax.inst[3] ;
 wire \minimax.inst[4] ;
 wire \minimax.inst[5] ;
 wire \minimax.inst[6] ;
 wire \minimax.inst[7] ;
 wire \minimax.inst[8] ;
 wire \minimax.inst[9] ;
 wire \minimax.inst_regce ;
 wire \minimax.microcode ;
 wire \minimax.op16_lw ;
 wire \minimax.op16_lwsp ;
 wire \minimax.op16_slli_setrd ;
 wire \minimax.op16_slli_setrs ;
 wire \minimax.pc_execute[1] ;
 wire \minimax.pc_execute[2] ;
 wire \minimax.pc_execute[3] ;
 wire \minimax.pc_execute[4] ;
 wire \minimax.pc_execute[5] ;
 wire \minimax.pc_execute[6] ;
 wire \minimax.pc_execute[7] ;
 wire \minimax.pc_execute[8] ;
 wire \minimax.pc_execute[9] ;
 wire \minimax.pc_fetch[1] ;
 wire \minimax.pc_fetch[2] ;
 wire \minimax.pc_fetch[3] ;
 wire \minimax.pc_fetch[4] ;
 wire \minimax.pc_fetch[5] ;
 wire \minimax.pc_fetch[6] ;
 wire \minimax.pc_fetch[7] ;
 wire \minimax.pc_fetch[8] ;
 wire \minimax.pc_fetch[9] ;
 wire \minimax.pc_fetch_dly[1] ;
 wire \minimax.pc_fetch_dly[2] ;
 wire \minimax.pc_fetch_dly[3] ;
 wire \minimax.pc_fetch_dly[4] ;
 wire \minimax.pc_fetch_dly[5] ;
 wire \minimax.pc_fetch_dly[6] ;
 wire \minimax.pc_fetch_dly[7] ;
 wire \minimax.pc_fetch_dly[8] ;
 wire \minimax.pc_fetch_dly[9] ;
 wire \minimax.regD_ex[0] ;
 wire \minimax.regD_ex[10] ;
 wire \minimax.regD_ex[11] ;
 wire \minimax.regD_ex[12] ;
 wire \minimax.regD_ex[13] ;
 wire \minimax.regD_ex[14] ;
 wire \minimax.regD_ex[15] ;
 wire \minimax.regD_ex[16] ;
 wire \minimax.regD_ex[17] ;
 wire \minimax.regD_ex[18] ;
 wire \minimax.regD_ex[19] ;
 wire \minimax.regD_ex[1] ;
 wire \minimax.regD_ex[20] ;
 wire \minimax.regD_ex[21] ;
 wire \minimax.regD_ex[22] ;
 wire \minimax.regD_ex[23] ;
 wire \minimax.regD_ex[24] ;
 wire \minimax.regD_ex[25] ;
 wire \minimax.regD_ex[26] ;
 wire \minimax.regD_ex[27] ;
 wire \minimax.regD_ex[28] ;
 wire \minimax.regD_ex[29] ;
 wire \minimax.regD_ex[2] ;
 wire \minimax.regD_ex[30] ;
 wire \minimax.regD_ex[31] ;
 wire \minimax.regD_ex[3] ;
 wire \minimax.regD_ex[4] ;
 wire \minimax.regD_ex[5] ;
 wire \minimax.regD_ex[6] ;
 wire \minimax.regD_ex[7] ;
 wire \minimax.regD_ex[8] ;
 wire \minimax.regD_ex[9] ;
 wire \minimax.regD_uc[0] ;
 wire \minimax.regD_uc[10] ;
 wire \minimax.regD_uc[11] ;
 wire \minimax.regD_uc[12] ;
 wire \minimax.regD_uc[13] ;
 wire \minimax.regD_uc[14] ;
 wire \minimax.regD_uc[15] ;
 wire \minimax.regD_uc[16] ;
 wire \minimax.regD_uc[17] ;
 wire \minimax.regD_uc[18] ;
 wire \minimax.regD_uc[19] ;
 wire \minimax.regD_uc[1] ;
 wire \minimax.regD_uc[20] ;
 wire \minimax.regD_uc[21] ;
 wire \minimax.regD_uc[22] ;
 wire \minimax.regD_uc[23] ;
 wire \minimax.regD_uc[24] ;
 wire \minimax.regD_uc[25] ;
 wire \minimax.regD_uc[26] ;
 wire \minimax.regD_uc[27] ;
 wire \minimax.regD_uc[28] ;
 wire \minimax.regD_uc[29] ;
 wire \minimax.regD_uc[2] ;
 wire \minimax.regD_uc[30] ;
 wire \minimax.regD_uc[31] ;
 wire \minimax.regD_uc[3] ;
 wire \minimax.regD_uc[4] ;
 wire \minimax.regD_uc[5] ;
 wire \minimax.regD_uc[6] ;
 wire \minimax.regD_uc[7] ;
 wire \minimax.regD_uc[8] ;
 wire \minimax.regD_uc[9] ;
 wire \minimax.regS_ex[0] ;
 wire \minimax.regS_ex[10] ;
 wire \minimax.regS_ex[11] ;
 wire \minimax.regS_ex[12] ;
 wire \minimax.regS_ex[13] ;
 wire \minimax.regS_ex[14] ;
 wire \minimax.regS_ex[15] ;
 wire \minimax.regS_ex[16] ;
 wire \minimax.regS_ex[17] ;
 wire \minimax.regS_ex[18] ;
 wire \minimax.regS_ex[19] ;
 wire \minimax.regS_ex[1] ;
 wire \minimax.regS_ex[20] ;
 wire \minimax.regS_ex[21] ;
 wire \minimax.regS_ex[22] ;
 wire \minimax.regS_ex[23] ;
 wire \minimax.regS_ex[24] ;
 wire \minimax.regS_ex[25] ;
 wire \minimax.regS_ex[26] ;
 wire \minimax.regS_ex[27] ;
 wire \minimax.regS_ex[28] ;
 wire \minimax.regS_ex[29] ;
 wire \minimax.regS_ex[2] ;
 wire \minimax.regS_ex[30] ;
 wire \minimax.regS_ex[31] ;
 wire \minimax.regS_ex[3] ;
 wire \minimax.regS_ex[4] ;
 wire \minimax.regS_ex[5] ;
 wire \minimax.regS_ex[6] ;
 wire \minimax.regS_ex[7] ;
 wire \minimax.regS_ex[8] ;
 wire \minimax.regS_ex[9] ;
 wire \minimax.regS_uc[0] ;
 wire \minimax.regS_uc[10] ;
 wire \minimax.regS_uc[11] ;
 wire \minimax.regS_uc[12] ;
 wire \minimax.regS_uc[13] ;
 wire \minimax.regS_uc[14] ;
 wire \minimax.regS_uc[15] ;
 wire \minimax.regS_uc[16] ;
 wire \minimax.regS_uc[17] ;
 wire \minimax.regS_uc[18] ;
 wire \minimax.regS_uc[19] ;
 wire \minimax.regS_uc[1] ;
 wire \minimax.regS_uc[20] ;
 wire \minimax.regS_uc[21] ;
 wire \minimax.regS_uc[22] ;
 wire \minimax.regS_uc[23] ;
 wire \minimax.regS_uc[24] ;
 wire \minimax.regS_uc[25] ;
 wire \minimax.regS_uc[26] ;
 wire \minimax.regS_uc[27] ;
 wire \minimax.regS_uc[28] ;
 wire \minimax.regS_uc[29] ;
 wire \minimax.regS_uc[2] ;
 wire \minimax.regS_uc[30] ;
 wire \minimax.regS_uc[31] ;
 wire \minimax.regS_uc[3] ;
 wire \minimax.regS_uc[4] ;
 wire \minimax.regS_uc[5] ;
 wire \minimax.regS_uc[6] ;
 wire \minimax.regS_uc[7] ;
 wire \minimax.regS_uc[8] ;
 wire \minimax.regS_uc[9] ;
 wire net360;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;

 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2157_ (.I(\minimax.inst[1] ),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2158_ (.I(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2159_ (.I(_1625_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2160_ (.I(\minimax.inst[13] ),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2161_ (.I(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2162_ (.I(_1628_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2163_ (.I(\minimax.inst[14] ),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2164_ (.I(_1630_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2165_ (.A1(_1629_),
    .A2(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2166_ (.A1(\minimax.inst[15] ),
    .A2(\minimax.inst[0] ),
    .A3(\minimax.bubble1 ),
    .A4(\minimax.bubble2 ),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2167_ (.A1(_1632_),
    .A2(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2168_ (.I(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2169_ (.A1(_1626_),
    .A2(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2170_ (.I(_1636_),
    .Z(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2171_ (.I(\minimax.inst[1] ),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2172_ (.I(_1637_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2173_ (.I(_1635_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2174_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_1638_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2176_ (.I(_1641_),
    .Z(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2177_ (.I(_1640_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2178_ (.I(\minimax.inst[3] ),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2179_ (.I(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2180_ (.I(\minimax.inst[2] ),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2181_ (.I(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2182_ (.I(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2183_ (.I(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2184_ (.I(\minimax.inst[12] ),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2185_ (.I(_1648_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2186_ (.I(_1649_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2187_ (.A1(\minimax.inst[13] ),
    .A2(\minimax.inst[14] ),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2188_ (.I(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _2189_ (.A1(\minimax.inst[4] ),
    .A2(\minimax.inst[5] ),
    .A3(\minimax.inst[6] ),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2190_ (.I(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2191_ (.A1(_1626_),
    .A2(_1652_),
    .A3(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2192_ (.A1(_1650_),
    .A2(_1633_),
    .A3(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2193_ (.A1(_1643_),
    .A2(_1647_),
    .A3(_1656_),
    .ZN(\minimax.op16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2194_ (.I(\minimax.inst[3] ),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2195_ (.I(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2196_ (.A1(_1658_),
    .A2(_1646_),
    .A3(_1656_),
    .ZN(\minimax.op16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2197_ (.A1(_1627_),
    .A2(\minimax.inst[14] ),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2198_ (.I(_1659_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _2199_ (.I(\minimax.inst[15] ),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2200_ (.I(\minimax.inst[0] ),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2201_ (.I(\minimax.bubble1 ),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _2202_ (.A1(_1624_),
    .A2(_1663_),
    .A3(\minimax.bubble2 ),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2203_ (.A1(_1661_),
    .A2(_1662_),
    .A3(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2204_ (.A1(_1660_),
    .A2(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2205_ (.I(\minimax.inst[12] ),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2206_ (.I(\minimax.inst[4] ),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2207_ (.I(\minimax.inst[5] ),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2208_ (.I(\minimax.inst[6] ),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2209_ (.A1(_1668_),
    .A2(_1669_),
    .A3(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2210_ (.A1(_1657_),
    .A2(_1644_),
    .A3(_1667_),
    .A4(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2211_ (.A1(_1669_),
    .A2(_1670_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2212_ (.A1(net410),
    .A2(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2213_ (.I(\minimax.inst[11] ),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2214_ (.I0(net376),
    .I1(_1674_),
    .S(_1675_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2215_ (.I(\minimax.inst[15] ),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2216_ (.I(\minimax.bubble2 ),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _2217_ (.A1(\minimax.inst[0] ),
    .A2(_1624_),
    .A3(_1663_),
    .A4(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2218_ (.A1(_1628_),
    .A2(_1630_),
    .A3(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2219_ (.I(_1675_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2220_ (.A1(net411),
    .A2(_1673_),
    .B(_1651_),
    .C(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2221_ (.A1(_1677_),
    .A2(_1651_),
    .A3(net383),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2222_ (.A1(_1677_),
    .A2(_1680_),
    .B1(_1682_),
    .B2(_1665_),
    .C(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2223_ (.A1(_1666_),
    .A2(_1676_),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2224_ (.I(_1685_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _2225_ (.I(\minimax.inst[8] ),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2226_ (.A1(\minimax.inst[7] ),
    .A2(\minimax.inst[9] ),
    .A3(net410),
    .A4(_1675_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2227_ (.A1(_1687_),
    .A2(net372),
    .A3(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2228_ (.I(\minimax.inst[15] ),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2229_ (.I(_1662_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2230_ (.A1(_1690_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2231_ (.A1(\minimax.inst[3] ),
    .A2(_1644_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2232_ (.A1(_1637_),
    .A2(\minimax.inst[12] ),
    .A3(_1660_),
    .A4(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2233_ (.A1(_1663_),
    .A2(_1678_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2234_ (.I(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2235_ (.A1(_1689_),
    .A2(_1692_),
    .A3(_1694_),
    .B(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2236_ (.I(_1667_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2237_ (.A1(_1624_),
    .A2(_1633_),
    .A3(_1659_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2238_ (.A1(_1657_),
    .A2(\minimax.inst[2] ),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2239_ (.A1(_1698_),
    .A2(_1653_),
    .A3(_1699_),
    .A4(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2240_ (.I(\minimax.inst[0] ),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2241_ (.A1(_1702_),
    .A2(_1625_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2242_ (.I(\minimax.inst[14] ),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2243_ (.A1(_1690_),
    .A2(_1704_),
    .B(_1627_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2244_ (.I(_1627_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2245_ (.A1(_1661_),
    .A2(_1637_),
    .B(_1706_),
    .C(\minimax.inst[14] ),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _2246_ (.A1(_1703_),
    .A2(_1705_),
    .B1(_1699_),
    .B2(_1672_),
    .C1(_1707_),
    .C2(_1702_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _2247_ (.A1(_1697_),
    .A2(_1701_),
    .A3(_1708_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2248_ (.A1(\minimax.inst[3] ),
    .A2(_1644_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2249_ (.A1(_1698_),
    .A2(_1654_),
    .A3(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2250_ (.A1(_1690_),
    .A2(_1662_),
    .A3(_1637_),
    .A4(_1695_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2251_ (.A1(_1624_),
    .A2(net398),
    .A3(net391),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2252_ (.A1(_1661_),
    .A2(_1702_),
    .A3(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2253_ (.A1(_1652_),
    .A2(_1711_),
    .A3(_1712_),
    .B1(_1714_),
    .B2(_1628_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2254_ (.A1(_1637_),
    .A2(_1659_),
    .A3(_1671_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2255_ (.I(\minimax.inst[8] ),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _2256_ (.A1(\minimax.inst[7] ),
    .A2(\minimax.inst[9] ),
    .A3(\minimax.inst[10] ),
    .A4(\minimax.inst[11] ),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2257_ (.A1(_1717_),
    .A2(_1667_),
    .A3(_1653_),
    .A4(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2258_ (.A1(_1690_),
    .A2(_1662_),
    .A3(_1695_),
    .A4(_1693_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2259_ (.A1(_1669_),
    .A2(net406),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2260_ (.A1(_1668_),
    .A2(\minimax.inst[12] ),
    .A3(_1721_),
    .A4(_1693_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _2261_ (.A1(_1716_),
    .A2(_1719_),
    .A3(_1720_),
    .B1(net408),
    .B2(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2262_ (.A1(_1715_),
    .A2(_1723_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2263_ (.I(\minimax.microcode ),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2264_ (.A1(_1725_),
    .A2(\minimax.dly16_slli_setrd ),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2265_ (.A1(_1686_),
    .A2(net380),
    .A3(_1724_),
    .B(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2266_ (.I(_1727_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2267_ (.I(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2268_ (.I(_1729_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2269_ (.I(_1730_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2270_ (.I(_1731_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2271_ (.I(_1732_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2272_ (.I0(\minimax.regD_ex[2] ),
    .I1(\minimax.regD_uc[2] ),
    .S(_1733_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2273_ (.I(_1734_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2274_ (.A1(\minimax.regD_uc[1] ),
    .A2(_1732_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2275_ (.A1(\minimax.microcode ),
    .A2(\minimax.dly16_slli_setrd ),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2276_ (.I(_1736_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2277_ (.I(_1686_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2278_ (.I(_1709_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2279_ (.I(_1724_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2280_ (.A1(_1738_),
    .A2(_1739_),
    .A3(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2281_ (.I(_1741_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2282_ (.A1(_1737_),
    .A2(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2283_ (.A1(\minimax.regD_ex[1] ),
    .A2(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2284_ (.A1(_1735_),
    .A2(_1744_),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2285_ (.I0(\minimax.regD_ex[0] ),
    .I1(\minimax.regD_uc[0] ),
    .S(_1733_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2286_ (.I(_1745_),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2287_ (.I(_1639_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2288_ (.A1(\minimax.pc_fetch[2] ),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2289_ (.I(_1634_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2290_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2291_ (.I(_1668_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2292_ (.I(_1664_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2293_ (.A1(_1691_),
    .A2(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2294_ (.I(net410),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2295_ (.A1(_1690_),
    .A2(_1627_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2296_ (.A1(_1753_),
    .A2(_1681_),
    .A3(_1651_),
    .B(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2297_ (.A1(_1752_),
    .A2(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2298_ (.I(_1756_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2299_ (.A1(_1750_),
    .A2(_1757_),
    .B(\minimax.regS_ex[2] ),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2300_ (.I(_1710_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2301_ (.A1(_1759_),
    .A2(_1756_),
    .B(\minimax.regS_ex[1] ),
    .C(\minimax.regS_ex[0] ),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2302_ (.I(_1669_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2303_ (.I(net407),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2304_ (.I(_1666_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2305_ (.I(_1753_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2306_ (.I(_1675_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2307_ (.A1(_1764_),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2308_ (.A1(_1761_),
    .A2(_1762_),
    .A3(_1763_),
    .A4(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2309_ (.A1(_1758_),
    .A2(_1760_),
    .A3(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2310_ (.I(_1661_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2311_ (.A1(_1769_),
    .A2(_1691_),
    .A3(_1652_),
    .A4(_1751_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2312_ (.I(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2313_ (.A1(_1753_),
    .A2(_1765_),
    .A3(_1721_),
    .A4(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2314_ (.I(_1668_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2315_ (.I(_1752_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2316_ (.I(_1755_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2317_ (.A1(_1774_),
    .A2(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2318_ (.I(\minimax.regS_uc[2] ),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2319_ (.A1(_1773_),
    .A2(_1776_),
    .B(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2320_ (.I(_1693_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2321_ (.A1(\minimax.regS_uc[1] ),
    .A2(\minimax.regS_uc[0] ),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2322_ (.A1(_1779_),
    .A2(_1776_),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2323_ (.A1(_1772_),
    .A2(_1778_),
    .A3(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2324_ (.A1(_1725_),
    .A2(\minimax.dly16_slli_setrs ),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2325_ (.A1(_1685_),
    .A2(_1709_),
    .A3(_1724_),
    .B(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2326_ (.I(net365),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2327_ (.I(_1785_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2328_ (.I0(_1768_),
    .I1(_1782_),
    .S(_1786_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(\minimax.regS_ex[1] ),
    .A2(\minimax.regS_ex[0] ),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2330_ (.A1(_1779_),
    .A2(_1776_),
    .B(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2331_ (.I(_1772_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2332_ (.A1(_1750_),
    .A2(_1757_),
    .B1(_1789_),
    .B2(_1790_),
    .C(\minimax.regS_ex[2] ),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2333_ (.A1(_1790_),
    .A2(_1781_),
    .B(_1778_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2334_ (.I0(_1791_),
    .I1(_1792_),
    .S(_1785_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2335_ (.A1(_1787_),
    .A2(_1793_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2336_ (.A1(_1628_),
    .A2(_1704_),
    .A3(_1717_),
    .A4(net369),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2337_ (.I(_1677_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2338_ (.A1(_1652_),
    .A2(_1795_),
    .B(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2339_ (.A1(_1682_),
    .A2(_1797_),
    .B(_1752_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2340_ (.A1(_1753_),
    .A2(_1675_),
    .A3(_1673_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2341_ (.A1(_1765_),
    .A2(net376),
    .B(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2342_ (.A1(_1654_),
    .A2(_1759_),
    .B(_1796_),
    .C(_1648_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2343_ (.A1(_1796_),
    .A2(net376),
    .B(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2344_ (.A1(_1691_),
    .A2(_1638_),
    .A3(_1696_),
    .A4(_1660_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2345_ (.A1(net379),
    .A2(_1800_),
    .B1(_1802_),
    .B2(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2346_ (.A1(_1798_),
    .A2(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2347_ (.I(_1726_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2348_ (.A1(\minimax.regD_uc[2] ),
    .A2(_1736_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2349_ (.A1(\minimax.regD_ex[2] ),
    .A2(_1806_),
    .B(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2350_ (.I(net384),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2351_ (.A1(_1809_),
    .A2(net368),
    .B(_1762_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2352_ (.I(_1750_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2353_ (.I(_1706_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2354_ (.A1(_1812_),
    .A2(_1704_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2355_ (.A1(_1813_),
    .A2(_1712_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2356_ (.I(\minimax.inst[9] ),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2357_ (.A1(_1811_),
    .A2(\minimax.op16_lwsp ),
    .B1(_1814_),
    .B2(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2358_ (.A1(_1805_),
    .A2(_1808_),
    .B(_1810_),
    .C(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2359_ (.A1(_1794_),
    .A2(_1817_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2360_ (.I(_1781_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2361_ (.I(_1785_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2362_ (.I0(_1760_),
    .I1(_1819_),
    .S(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2363_ (.I(\minimax.regD_uc[1] ),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2364_ (.A1(\minimax.regD_ex[1] ),
    .A2(_1806_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2365_ (.A1(\minimax.regD_ex[1] ),
    .A2(_1737_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _2366_ (.A1(_1677_),
    .A2(_1651_),
    .A3(_1679_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2367_ (.A1(_1769_),
    .A2(_1813_),
    .A3(net383),
    .B(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2368_ (.A1(net379),
    .A2(_1800_),
    .B1(_1682_),
    .B2(_1665_),
    .C(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2369_ (.A1(net378),
    .A2(net364),
    .A3(_1708_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2370_ (.A1(_1715_),
    .A2(_1723_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2371_ (.A1(_1827_),
    .A2(_1828_),
    .A3(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2372_ (.I(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2373_ (.I(_1805_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2374_ (.A1(_1822_),
    .A2(_1823_),
    .B1(_1824_),
    .B2(_1831_),
    .C(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2375_ (.A1(_1821_),
    .A2(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2376_ (.I(net374),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2377_ (.I(_1829_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_4 _2378_ (.A1(\minimax.microcode ),
    .A2(\minimax.dly16_slli_setrs ),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2379_ (.A1(_1644_),
    .A2(_1774_),
    .A3(_1775_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2380_ (.A1(\minimax.regS_ex[0] ),
    .A2(_1837_),
    .A3(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2381_ (.A1(_1835_),
    .A2(_1836_),
    .B(_1839_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2382_ (.I(net404),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2383_ (.A1(\minimax.regS_uc[0] ),
    .A2(_1838_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2384_ (.A1(_1835_),
    .A2(_1841_),
    .A3(_1836_),
    .A4(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2385_ (.I(_1783_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2386_ (.A1(\minimax.regS_uc[0] ),
    .A2(_1844_),
    .A3(_1838_),
    .B1(_1839_),
    .B2(_1841_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2387_ (.A1(_1840_),
    .A2(_1843_),
    .A3(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _2388_ (.I(_1704_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2389_ (.I(_1681_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2390_ (.I(_1677_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2391_ (.A1(_1847_),
    .A2(_1764_),
    .A3(_1848_),
    .B(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2392_ (.I(_1662_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2393_ (.A1(_1851_),
    .A2(_1629_),
    .A3(_1658_),
    .A4(net389),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2394_ (.A1(_1850_),
    .A2(_1852_),
    .B(_1837_),
    .C(\minimax.regS_ex[1] ),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2395_ (.A1(_1790_),
    .A2(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2396_ (.A1(_1738_),
    .A2(_1739_),
    .A3(_1740_),
    .B(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2397_ (.I(_1835_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2398_ (.I(_1841_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2399_ (.I(_1836_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2400_ (.A1(_1850_),
    .A2(_1852_),
    .B(\minimax.regS_uc[1] ),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2401_ (.A1(_1856_),
    .A2(_1857_),
    .A3(_1858_),
    .A4(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2402_ (.I(_1837_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2403_ (.I0(\minimax.regS_uc[1] ),
    .I1(_1859_),
    .S(_1790_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2404_ (.I(\minimax.regS_ex[1] ),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2405_ (.A1(_1658_),
    .A2(_1776_),
    .B1(_1861_),
    .B2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2406_ (.A1(_1861_),
    .A2(_1862_),
    .B1(_1864_),
    .B2(_1767_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2407_ (.A1(_1855_),
    .A2(_1860_),
    .A3(_1865_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2408_ (.A1(_1846_),
    .A2(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2409_ (.I(_1806_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2410_ (.A1(\minimax.regD_ex[0] ),
    .A2(_1868_),
    .B1(_1728_),
    .B2(\minimax.regD_uc[0] ),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2411_ (.A1(_1832_),
    .A2(_1869_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2412_ (.A1(_1840_),
    .A2(_1843_),
    .A3(_1845_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2413_ (.A1(_1821_),
    .A2(_1833_),
    .B1(_1871_),
    .B2(_1866_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2414_ (.A1(_1834_),
    .A2(_1867_),
    .B1(_1870_),
    .B2(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2415_ (.A1(_1818_),
    .A2(_1873_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_1749_),
    .A2(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2417_ (.I(net160),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2418_ (.I(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2419_ (.A1(_1747_),
    .A2(_1875_),
    .B(_1877_),
    .ZN(\bank1.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2420_ (.I0(\minimax.regD_ex[3] ),
    .I1(\minimax.regD_uc[3] ),
    .S(_1732_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2421_ (.I(_1878_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2422_ (.A1(\minimax.pc_fetch[3] ),
    .A2(_1746_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2423_ (.I(_1640_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2424_ (.I(_1817_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2425_ (.A1(_1834_),
    .A2(_1867_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2426_ (.A1(_1870_),
    .A2(_1872_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2427_ (.A1(_1882_),
    .A2(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2428_ (.A1(_1794_),
    .A2(_1817_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2429_ (.A1(_1884_),
    .A2(_1885_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2430_ (.A1(_1794_),
    .A2(_1881_),
    .B(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2431_ (.I(_1764_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2432_ (.A1(net367),
    .A2(_1814_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2433_ (.I0(\minimax.regD_ex[3] ),
    .I1(\minimax.regD_uc[3] ),
    .S(_1736_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2434_ (.I(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2435_ (.I(_1761_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2436_ (.A1(_1636_),
    .A2(net385),
    .B(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2437_ (.A1(_1888_),
    .A2(_1889_),
    .B1(_1891_),
    .B2(_1805_),
    .C(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2438_ (.I(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2439_ (.A1(_1761_),
    .A2(_1756_),
    .B(_1837_),
    .C(\minimax.regS_ex[3] ),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2440_ (.A1(_1686_),
    .A2(_1740_),
    .B(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2441_ (.A1(_1892_),
    .A2(_1757_),
    .B(\minimax.regS_uc[3] ),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2442_ (.A1(_1835_),
    .A2(_1841_),
    .A3(_1836_),
    .A4(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2443_ (.A1(_1892_),
    .A2(_1756_),
    .B(_1844_),
    .C(\minimax.regS_uc[3] ),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2444_ (.A1(_1739_),
    .A2(_1896_),
    .B(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2445_ (.A1(_1897_),
    .A2(_1899_),
    .A3(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2446_ (.A1(_1750_),
    .A2(_1759_),
    .B(_1757_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2447_ (.A1(\minimax.regS_ex[2] ),
    .A2(\minimax.regS_ex[1] ),
    .A3(\minimax.regS_ex[0] ),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2448_ (.A1(_1903_),
    .A2(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2449_ (.A1(\minimax.regS_uc[2] ),
    .A2(\minimax.regS_uc[1] ),
    .A3(\minimax.regS_uc[0] ),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2450_ (.A1(_1785_),
    .A2(_1903_),
    .A3(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2451_ (.I(_1772_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2452_ (.A1(_1786_),
    .A2(_1905_),
    .B(_1907_),
    .C(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2453_ (.A1(_1902_),
    .A2(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2454_ (.I(_1910_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2455_ (.A1(_1887_),
    .A2(_1895_),
    .A3(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2456_ (.A1(_1880_),
    .A2(_1912_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2457_ (.A1(_1879_),
    .A2(_1913_),
    .B(_1877_),
    .ZN(\bank1.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2458_ (.A1(_1794_),
    .A2(_1817_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2459_ (.A1(_1894_),
    .A2(_1902_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2460_ (.I0(_1787_),
    .I1(_1793_),
    .S(_1915_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2461_ (.A1(_1881_),
    .A2(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2462_ (.A1(_1914_),
    .A2(_1884_),
    .B(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2463_ (.A1(_1911_),
    .A2(_1918_),
    .B(_1895_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2464_ (.I(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2465_ (.A1(_1911_),
    .A2(_1918_),
    .B(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2466_ (.A1(_1796_),
    .A2(_1638_),
    .A3(_1847_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2467_ (.A1(_1769_),
    .A2(_1625_),
    .A3(_1631_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2468_ (.A1(_1691_),
    .A2(_1696_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2469_ (.A1(_1922_),
    .A2(_1923_),
    .B(_1629_),
    .C(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2470_ (.A1(_1680_),
    .A2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2471_ (.I(_1926_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2472_ (.A1(_1762_),
    .A2(_1636_),
    .B1(_1927_),
    .B2(_1765_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2473_ (.A1(_1798_),
    .A2(_1804_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2474_ (.I(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2475_ (.A1(\minimax.regD_ex[4] ),
    .A2(_1806_),
    .A3(_1930_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2476_ (.A1(\minimax.regD_uc[4] ),
    .A2(_1727_),
    .A3(_1929_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2477_ (.A1(_1928_),
    .A2(_1931_),
    .A3(_1932_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2478_ (.A1(\minimax.regS_ex[4] ),
    .A2(_1783_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2479_ (.A1(_1769_),
    .A2(_1753_),
    .A3(_1848_),
    .A4(_1652_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2480_ (.A1(_1628_),
    .A2(_1704_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2481_ (.A1(_1796_),
    .A2(_1687_),
    .A3(net397),
    .A4(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2482_ (.A1(_1935_),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _2483_ (.I(net406),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2484_ (.A1(_1702_),
    .A2(net401),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2485_ (.A1(_1754_),
    .A2(_1938_),
    .B(_1939_),
    .C(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2486_ (.A1(\minimax.regS_uc[4] ),
    .A2(net365),
    .B1(_1934_),
    .B2(_1830_),
    .C(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2487_ (.A1(_1668_),
    .A2(_1669_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2488_ (.A1(_1943_),
    .A2(_1779_),
    .B(net389),
    .C(_1851_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2489_ (.I(\minimax.regS_uc[3] ),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2490_ (.A1(_1945_),
    .A2(_1906_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2491_ (.A1(_1775_),
    .A2(_1944_),
    .B(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2492_ (.A1(_1837_),
    .A2(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2493_ (.A1(net377),
    .A2(_1828_),
    .A3(_1829_),
    .A4(_1947_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2494_ (.I(_1783_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2495_ (.I(\minimax.regS_ex[3] ),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2496_ (.A1(_1951_),
    .A2(_1904_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2497_ (.A1(_1775_),
    .A2(_1944_),
    .B(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2498_ (.A1(_1950_),
    .A2(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2499_ (.A1(_1686_),
    .A2(_1709_),
    .A3(_1724_),
    .B(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2500_ (.A1(_1790_),
    .A2(_1948_),
    .A3(_1949_),
    .A4(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2501_ (.A1(net405),
    .A2(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _2502_ (.A1(_1933_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2503_ (.A1(_1921_),
    .A2(_1958_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2504_ (.A1(\minimax.pc_fetch[4] ),
    .A2(_1748_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2505_ (.I(_1876_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2506_ (.A1(_1749_),
    .A2(_1959_),
    .B(_1960_),
    .C(_1961_),
    .ZN(\bank1.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2507_ (.A1(\minimax.pc_fetch[5] ),
    .A2(_1880_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2508_ (.A1(_1626_),
    .A2(_1635_),
    .B(_1926_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2509_ (.I0(\minimax.regD_ex[5] ),
    .I1(\minimax.regD_uc[5] ),
    .S(_1736_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2510_ (.A1(_1649_),
    .A2(_1963_),
    .B1(_1964_),
    .B2(_1929_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2511_ (.I(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2512_ (.A1(_1948_),
    .A2(_1949_),
    .A3(_1955_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2513_ (.A1(_1942_),
    .A2(_1967_),
    .B(_1767_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2514_ (.A1(_1648_),
    .A2(_1774_),
    .A3(_1755_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2515_ (.A1(net394),
    .A2(_1795_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2516_ (.A1(_1645_),
    .A2(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2517_ (.A1(\minimax.regS_ex[5] ),
    .A2(_1783_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2518_ (.A1(\minimax.regS_uc[5] ),
    .A2(_1785_),
    .B1(_1972_),
    .B2(_1830_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2519_ (.A1(_1969_),
    .A2(_1971_),
    .A3(_1973_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2520_ (.A1(_1966_),
    .A2(_1968_),
    .A3(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2521_ (.I(_1933_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2522_ (.I(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2523_ (.A1(_1977_),
    .A2(_1957_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2524_ (.A1(_1977_),
    .A2(_1957_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2525_ (.A1(_1921_),
    .A2(_1978_),
    .B(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2526_ (.A1(_1975_),
    .A2(_1980_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2527_ (.A1(_1749_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2528_ (.A1(_1962_),
    .A2(_1982_),
    .B(_1877_),
    .ZN(\bank1.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2529_ (.A1(\minimax.pc_fetch[6] ),
    .A2(_1880_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2530_ (.I(_1748_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2531_ (.A1(_1976_),
    .A2(_1957_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2532_ (.A1(_1895_),
    .A2(_1911_),
    .A3(_1975_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2533_ (.A1(_1968_),
    .A2(_1974_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2534_ (.A1(_1966_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2535_ (.A1(_1985_),
    .A2(_1986_),
    .B(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2536_ (.A1(_1818_),
    .A2(_1873_),
    .B1(_1916_),
    .B2(_1817_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2537_ (.A1(_1895_),
    .A2(_1911_),
    .B(_1958_),
    .C(_1975_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2538_ (.I(_1942_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2539_ (.A1(_1992_),
    .A2(_1956_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2540_ (.I(_1974_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2541_ (.A1(_1966_),
    .A2(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2542_ (.A1(_1965_),
    .A2(_1994_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2543_ (.A1(_1992_),
    .A2(_1956_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2544_ (.A1(_1993_),
    .A2(_1995_),
    .B1(_1996_),
    .B2(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2545_ (.A1(_1933_),
    .A2(_1957_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2546_ (.A1(_1894_),
    .A2(_1910_),
    .A3(_1999_),
    .A4(_1975_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2547_ (.A1(_1990_),
    .A2(_1991_),
    .B1(_1998_),
    .B2(_1976_),
    .C(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2548_ (.A1(_1989_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2549_ (.A1(_1645_),
    .A2(\minimax.op16_lwsp ),
    .B1(net367),
    .B2(_1892_),
    .C1(_1925_),
    .C2(\minimax.inst[7] ),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2550_ (.A1(\minimax.regD_uc[6] ),
    .A2(_1728_),
    .A3(_1930_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2551_ (.A1(\minimax.regD_ex[6] ),
    .A2(_1806_),
    .A3(_1930_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _2552_ (.A1(_2003_),
    .A2(_2004_),
    .A3(_2005_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2553_ (.I(_1992_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2554_ (.A1(_2007_),
    .A2(_1967_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _2555_ (.A1(_1971_),
    .A2(_1973_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2556_ (.I(_1969_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2557_ (.A1(_1761_),
    .A2(net400),
    .B(\minimax.regS_ex[6] ),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2558_ (.A1(_1761_),
    .A2(net400),
    .B(\minimax.regS_uc[6] ),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _2559_ (.I0(_2011_),
    .I1(_2012_),
    .S(net366),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2560_ (.A1(_2010_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2561_ (.I(_2014_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2562_ (.I(_1767_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2563_ (.I(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2564_ (.A1(_2008_),
    .A2(_2009_),
    .B(_2015_),
    .C(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2565_ (.I(_1908_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2566_ (.A1(_1950_),
    .A2(_1969_),
    .A3(_1953_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2567_ (.A1(_1686_),
    .A2(_1724_),
    .B(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2568_ (.A1(_1648_),
    .A2(_1752_),
    .A3(_1755_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2569_ (.A1(_1950_),
    .A2(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2570_ (.A1(_1709_),
    .A2(_2020_),
    .B1(_2023_),
    .B2(_1947_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2571_ (.A1(_1949_),
    .A2(_2021_),
    .A3(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2572_ (.A1(_1992_),
    .A2(_1971_),
    .A3(_1973_),
    .A4(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2573_ (.I(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2574_ (.A1(_2019_),
    .A2(_2027_),
    .B(net388),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2575_ (.A1(_2018_),
    .A2(_2028_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2576_ (.A1(_2006_),
    .A2(_2029_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2577_ (.A1(_2002_),
    .A2(_2030_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2578_ (.A1(_1984_),
    .A2(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2579_ (.I(_1876_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2580_ (.A1(_1983_),
    .A2(_2032_),
    .B(_2033_),
    .ZN(\bank1.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2581_ (.I(_1733_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _2582_ (.I0(\minimax.regD_ex[7] ),
    .I1(\minimax.regD_uc[7] ),
    .S(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2583_ (.I(_2035_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2584_ (.A1(\minimax.pc_fetch[7] ),
    .A2(_1880_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2585_ (.A1(_2003_),
    .A2(_2004_),
    .A3(_2005_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2586_ (.A1(_2002_),
    .A2(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2587_ (.A1(_2029_),
    .A2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2588_ (.A1(_2002_),
    .A2(_2037_),
    .B(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2589_ (.I(_1930_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2590_ (.A1(\minimax.regD_ex[7] ),
    .A2(_1868_),
    .A3(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2591_ (.I(_1717_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2592_ (.A1(_1642_),
    .A2(\minimax.op16_lwsp ),
    .B1(_1925_),
    .B2(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2593_ (.A1(\minimax.regD_uc[7] ),
    .A2(_1728_),
    .A3(_1930_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _2594_ (.A1(_2042_),
    .A2(_2044_),
    .A3(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2595_ (.I(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2596_ (.A1(_1992_),
    .A2(_1971_),
    .A3(_1973_),
    .A4(_2025_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2597_ (.I(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2598_ (.I(_2049_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2599_ (.A1(net388),
    .A2(_2050_),
    .B(_2017_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2600_ (.I(\minimax.regS_ex[7] ),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2601_ (.A1(_1849_),
    .A2(_1851_),
    .A3(net389),
    .A4(_1936_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2602_ (.A1(_1717_),
    .A2(\minimax.inst[3] ),
    .A3(net370),
    .A4(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2603_ (.A1(_2052_),
    .A2(_1950_),
    .A3(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2604_ (.A1(_1835_),
    .A2(_1836_),
    .B(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2605_ (.A1(_1642_),
    .A2(_1970_),
    .B(\minimax.regS_uc[7] ),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2606_ (.A1(net371),
    .A2(net390),
    .A3(_1829_),
    .A4(_2057_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2607_ (.I(_2054_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2608_ (.A1(\minimax.regS_uc[7] ),
    .A2(_1950_),
    .A3(_2059_),
    .B1(_2055_),
    .B2(_1841_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2609_ (.A1(_2056_),
    .A2(_2058_),
    .A3(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2610_ (.A1(_2010_),
    .A2(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2611_ (.A1(_2051_),
    .A2(_2062_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2612_ (.A1(_2040_),
    .A2(_2047_),
    .A3(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2613_ (.A1(_1984_),
    .A2(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2614_ (.A1(_2036_),
    .A2(_2065_),
    .B(_2033_),
    .ZN(\bank1.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _2615_ (.I0(\minimax.regD_ex[8] ),
    .I1(\minimax.regD_uc[8] ),
    .S(_2034_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2616_ (.I(_2066_),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2617_ (.A1(\minimax.pc_fetch[8] ),
    .A2(_1880_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _2618_ (.I(_1815_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2619_ (.A1(\minimax.regD_uc[8] ),
    .A2(_1737_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2620_ (.A1(\minimax.regD_ex[8] ),
    .A2(_1868_),
    .B(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2621_ (.A1(_2068_),
    .A2(net386),
    .B1(_1832_),
    .B2(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2622_ (.I(_1786_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2623_ (.A1(\minimax.regS_uc[8] ),
    .A2(_2072_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2624_ (.A1(_2043_),
    .A2(net370),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2625_ (.A1(net395),
    .A2(_0075_),
    .A3(_1936_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _2626_ (.I(\minimax.regS_ex[8] ),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2627_ (.A1(_0077_),
    .A2(_1861_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2628_ (.A1(_1811_),
    .A2(_0076_),
    .B1(_0078_),
    .B2(_1831_),
    .C(_2022_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2629_ (.A1(_0074_),
    .A2(_0079_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2630_ (.A1(_1642_),
    .A2(net400),
    .B(\minimax.regS_ex[7] ),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2631_ (.A1(_2011_),
    .A2(_0081_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2632_ (.A1(_2012_),
    .A2(_2057_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2633_ (.I(_2072_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _2634_ (.I0(_0082_),
    .I1(_0083_),
    .S(_0084_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2635_ (.A1(_2007_),
    .A2(_2025_),
    .A3(_0085_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2636_ (.A1(_2011_),
    .A2(_0081_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2637_ (.A1(_2012_),
    .A2(_2057_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2638_ (.I0(_0087_),
    .I1(_0088_),
    .S(_1820_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2639_ (.I(_0074_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2640_ (.I(_0079_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2641_ (.A1(_2071_),
    .A2(_0089_),
    .A3(_0090_),
    .A4(_0091_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2642_ (.A1(_2071_),
    .A2(_0080_),
    .A3(_0086_),
    .B(_0092_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2643_ (.A1(_2071_),
    .A2(_0080_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2644_ (.I0(_0093_),
    .I1(_0094_),
    .S(_2017_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2645_ (.A1(\minimax.regS_uc[8] ),
    .A2(_1820_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2646_ (.A1(_1811_),
    .A2(_0076_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2647_ (.A1(_0077_),
    .A2(_1820_),
    .B(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2648_ (.A1(_0096_),
    .A2(_0098_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2649_ (.A1(_2050_),
    .A2(_0085_),
    .A3(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2650_ (.I(_2019_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2651_ (.I(_2027_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2652_ (.I(_0080_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2653_ (.A1(_0101_),
    .A2(_0102_),
    .A3(_0103_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2654_ (.I(_2070_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2655_ (.A1(_1815_),
    .A2(_1809_),
    .B1(_2041_),
    .B2(_0105_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2656_ (.I(_0106_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2657_ (.A1(_0100_),
    .A2(_0104_),
    .B(_0107_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2658_ (.A1(_1763_),
    .A2(_1766_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2659_ (.A1(_1721_),
    .A2(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(_0110_),
    .A2(_0106_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2661_ (.A1(_2009_),
    .A2(_0107_),
    .A3(_0103_),
    .A4(_0086_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2662_ (.A1(_2009_),
    .A2(_0103_),
    .A3(_0111_),
    .B(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2663_ (.A1(_0095_),
    .A2(_0108_),
    .A3(_0113_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2664_ (.A1(_2042_),
    .A2(_2044_),
    .A3(_2045_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2665_ (.A1(_0115_),
    .A2(_2063_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2666_ (.A1(_0115_),
    .A2(_2063_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2667_ (.A1(_2040_),
    .A2(_0116_),
    .B(_0117_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2668_ (.A1(_0114_),
    .A2(_0118_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(_1984_),
    .A2(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2670_ (.A1(_2067_),
    .A2(_0120_),
    .B(_2033_),
    .ZN(\bank1.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _2671_ (.I0(\minimax.regD_ex[9] ),
    .I1(\minimax.regD_uc[9] ),
    .S(_2034_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2672_ (.I(_0121_),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2673_ (.A1(_2010_),
    .A2(_2013_),
    .A3(_2061_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2674_ (.A1(_2026_),
    .A2(_0099_),
    .A3(_0122_),
    .B(_2019_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2675_ (.A1(\minimax.regS_ex[9] ),
    .A2(_1844_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2676_ (.I(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2677_ (.A1(_1849_),
    .A2(_1631_),
    .A3(_1687_),
    .A4(net397),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2678_ (.A1(_1775_),
    .A2(_0126_),
    .B(_1648_),
    .C(_1774_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _2679_ (.I(_0127_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2680_ (.A1(\minimax.regS_uc[9] ),
    .A2(_1820_),
    .B1(_0125_),
    .B2(_1831_),
    .C(_0128_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2681_ (.I(_1764_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2682_ (.A1(\minimax.regD_uc[9] ),
    .A2(_1737_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2683_ (.A1(\minimax.regD_ex[9] ),
    .A2(_1868_),
    .B(_0131_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2684_ (.A1(_1798_),
    .A2(_1804_),
    .B(_0132_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2685_ (.A1(_0130_),
    .A2(_1809_),
    .B(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2686_ (.A1(_0123_),
    .A2(net409),
    .A3(_0134_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2687_ (.A1(_2056_),
    .A2(_2058_),
    .A3(_2060_),
    .B(_2010_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2688_ (.A1(_2016_),
    .A2(_0136_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2689_ (.A1(_2015_),
    .A2(_0137_),
    .B(_2046_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2690_ (.I(_2011_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2691_ (.I(_2012_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2692_ (.I0(_0139_),
    .I1(_0140_),
    .S(_1786_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2693_ (.A1(_2022_),
    .A2(_0141_),
    .B(_1908_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2694_ (.A1(_2006_),
    .A2(_2014_),
    .B1(_2048_),
    .B2(_2016_),
    .C(_0142_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2695_ (.A1(_2037_),
    .A2(_0138_),
    .B1(_0143_),
    .B2(_2062_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2696_ (.A1(_0141_),
    .A2(_2026_),
    .B(_1908_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2697_ (.I(_0136_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2698_ (.A1(_2014_),
    .A2(_2026_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2699_ (.A1(_1908_),
    .A2(_0136_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2700_ (.A1(_2010_),
    .A2(_2013_),
    .B(_2048_),
    .C(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2701_ (.A1(_2022_),
    .A2(_0141_),
    .A3(_0136_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _2702_ (.A1(_0145_),
    .A2(_0146_),
    .A3(_0147_),
    .B1(_0149_),
    .B2(_0150_),
    .B3(_0115_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2703_ (.A1(_1985_),
    .A2(_1986_),
    .B1(_0144_),
    .B2(_0151_),
    .C(_1988_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2704_ (.A1(_2001_),
    .A2(_0152_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2705_ (.I(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2706_ (.A1(_2051_),
    .A2(_0146_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2707_ (.A1(_2018_),
    .A2(_2028_),
    .B1(_2047_),
    .B2(_0101_),
    .C(_2006_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2708_ (.A1(_0145_),
    .A2(_2062_),
    .B(_2047_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2709_ (.A1(_2018_),
    .A2(_2028_),
    .B1(_2046_),
    .B2(_0148_),
    .C(_2006_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2710_ (.A1(_0155_),
    .A2(_0156_),
    .B1(_0157_),
    .B2(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2711_ (.A1(_0114_),
    .A2(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2712_ (.A1(_0090_),
    .A2(_0091_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2713_ (.I(_0161_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2714_ (.I(_0101_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2715_ (.I(_0163_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2716_ (.I(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2717_ (.I(_0165_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2718_ (.A1(_2050_),
    .A2(_0085_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2719_ (.A1(_0166_),
    .A2(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2720_ (.A1(_0162_),
    .A2(_0168_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2721_ (.I(_2071_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2722_ (.A1(_0154_),
    .A2(_0160_),
    .B1(_0169_),
    .B2(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2723_ (.A1(_0135_),
    .A2(_0171_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2724_ (.A1(\minimax.pc_fetch[9] ),
    .A2(_1748_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2725_ (.A1(_1749_),
    .A2(_0172_),
    .B(_0173_),
    .C(_1961_),
    .ZN(\bank1.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2726_ (.I0(\minimax.regD_ex[10] ),
    .I1(\minimax.regD_uc[10] ),
    .S(_1727_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2727_ (.I(_0174_),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2728_ (.A1(_2041_),
    .A2(net3),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2729_ (.A1(_0074_),
    .A2(_0079_),
    .A3(_0129_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2730_ (.A1(_2026_),
    .A2(_0089_),
    .A3(_0176_),
    .B(_2019_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2731_ (.I(_1861_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2732_ (.A1(_1741_),
    .A2(_0178_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2733_ (.A1(\minimax.regS_uc[10] ),
    .A2(_0084_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2734_ (.A1(\minimax.regS_ex[10] ),
    .A2(_0179_),
    .B(_0128_),
    .C(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _2735_ (.A1(_0175_),
    .A2(_0177_),
    .A3(_0181_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2736_ (.A1(_0095_),
    .A2(_0108_),
    .A3(_0113_),
    .B(_0135_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2737_ (.A1(_0159_),
    .A2(_0183_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2738_ (.I(_0129_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2739_ (.A1(_0103_),
    .A2(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2740_ (.I(_0127_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2741_ (.I(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2742_ (.I(_2072_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2743_ (.I(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2744_ (.I(_1831_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2745_ (.A1(\minimax.regS_uc[9] ),
    .A2(_0190_),
    .B1(_0125_),
    .B2(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2746_ (.A1(_0188_),
    .A2(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2747_ (.A1(_0193_),
    .A2(_0134_),
    .B(_0107_),
    .C(_0161_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2748_ (.I(_1888_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2749_ (.A1(_0195_),
    .A2(net387),
    .B1(_1832_),
    .B2(_0132_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2750_ (.A1(_0129_),
    .A2(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2751_ (.A1(_0090_),
    .A2(_0091_),
    .B(_0134_),
    .C(_2016_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2752_ (.A1(_0197_),
    .A2(_0198_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2753_ (.A1(_0123_),
    .A2(_0186_),
    .B1(_0194_),
    .B2(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2754_ (.A1(_0185_),
    .A2(_0134_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2755_ (.A1(_0185_),
    .A2(_0134_),
    .B(_0107_),
    .C(_0103_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2756_ (.I(_2019_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2757_ (.A1(_0201_),
    .A2(_0202_),
    .B(_0203_),
    .C(_0167_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2758_ (.A1(_0200_),
    .A2(_0204_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2759_ (.A1(_0154_),
    .A2(_0184_),
    .B(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2760_ (.A1(_0182_),
    .A2(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2761_ (.A1(net160),
    .A2(_1639_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2762_ (.I(_0208_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2763_ (.A1(_0207_),
    .A2(_0209_),
    .ZN(\bank1.addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2764_ (.I0(\minimax.regD_ex[11] ),
    .I1(\minimax.regD_uc[11] ),
    .S(_1727_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2765_ (.I(_0210_),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2766_ (.I0(\minimax.regD_ex[12] ),
    .I1(\minimax.regD_uc[12] ),
    .S(_1729_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2767_ (.I(_0211_),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2768_ (.A1(_2041_),
    .A2(net4),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2769_ (.I(_0212_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2770_ (.I(\minimax.regS_ex[11] ),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2771_ (.I(\minimax.regS_uc[11] ),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2772_ (.I0(_0214_),
    .I1(_0215_),
    .S(_2072_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2773_ (.A1(_0188_),
    .A2(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2774_ (.I(_0122_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2775_ (.I(_1844_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2776_ (.A1(\minimax.regS_ex[9] ),
    .A2(\minimax.regS_ex[10] ),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2777_ (.A1(_0219_),
    .A2(_0187_),
    .A3(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2778_ (.A1(_1856_),
    .A2(_1858_),
    .B(_0221_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2779_ (.A1(\minimax.regS_uc[9] ),
    .A2(\minimax.regS_uc[10] ),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(_0127_),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2781_ (.A1(_1738_),
    .A2(_1739_),
    .A3(_1740_),
    .A4(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2782_ (.A1(_1861_),
    .A2(_0187_),
    .A3(_0223_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2783_ (.A1(_1857_),
    .A2(_0221_),
    .B(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2784_ (.A1(_0222_),
    .A2(_0225_),
    .A3(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _2785_ (.A1(_0096_),
    .A2(_0098_),
    .A3(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2786_ (.A1(_2027_),
    .A2(_0218_),
    .A3(_0229_),
    .B(_0101_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2787_ (.A1(_0213_),
    .A2(_0217_),
    .A3(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2788_ (.I(_1892_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2789_ (.I(_1762_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2790_ (.I(_1765_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2791_ (.A1(_1764_),
    .A2(_0234_),
    .A3(_1771_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2792_ (.A1(_0232_),
    .A2(_0233_),
    .A3(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2793_ (.A1(_0236_),
    .A2(_0217_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2794_ (.I(_2041_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2795_ (.A1(_0238_),
    .A2(net4),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2796_ (.I0(\minimax.regS_ex[11] ),
    .I1(\minimax.regS_uc[11] ),
    .S(_0084_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2797_ (.A1(_0239_),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2798_ (.I(_0150_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2799_ (.A1(_0096_),
    .A2(_0098_),
    .A3(_0228_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2800_ (.I(_0243_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2801_ (.A1(_2050_),
    .A2(_0242_),
    .A3(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _2802_ (.A1(_0213_),
    .A2(_0237_),
    .B1(_0241_),
    .B2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2803_ (.A1(_2016_),
    .A2(_0128_),
    .A3(_0240_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2804_ (.A1(_2027_),
    .A2(_0218_),
    .A3(_0229_),
    .B(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2805_ (.A1(_2049_),
    .A2(_0150_),
    .A3(_0243_),
    .A4(_0240_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2806_ (.A1(_0212_),
    .A2(_0248_),
    .A3(_0249_),
    .A4(_0237_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2807_ (.A1(_0231_),
    .A2(_0246_),
    .A3(_0250_),
    .B(_0182_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2808_ (.A1(_0159_),
    .A2(_0183_),
    .A3(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2809_ (.A1(_0153_),
    .A2(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2810_ (.I(_0175_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2811_ (.A1(_0254_),
    .A2(_0181_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2812_ (.I(\minimax.regS_ex[10] ),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _2813_ (.I(_2072_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2814_ (.A1(\minimax.regS_uc[10] ),
    .A2(_0189_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2815_ (.A1(_0256_),
    .A2(_0257_),
    .B(_0188_),
    .C(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(_0175_),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2817_ (.I0(_0255_),
    .I1(_0260_),
    .S(_0177_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2818_ (.A1(_0177_),
    .A2(_0181_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2819_ (.A1(_0254_),
    .A2(_0262_),
    .B1(_0200_),
    .B2(_0204_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2820_ (.A1(_0248_),
    .A2(_0249_),
    .A3(_0237_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2821_ (.A1(_0213_),
    .A2(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2822_ (.A1(_0261_),
    .A2(_0263_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2823_ (.I(_0239_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2824_ (.A1(_0248_),
    .A2(_0249_),
    .A3(_0237_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2825_ (.A1(_0267_),
    .A2(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2826_ (.A1(_0266_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2827_ (.I(_0238_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2828_ (.I(_0216_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2829_ (.A1(_2049_),
    .A2(_0150_),
    .A3(_0244_),
    .A4(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2830_ (.I(\minimax.regS_ex[12] ),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2831_ (.A1(_1645_),
    .A2(_0075_),
    .A3(_2053_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2832_ (.A1(_0274_),
    .A2(_0219_),
    .A3(_0127_),
    .A4(_0275_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2833_ (.A1(_1738_),
    .A2(_1740_),
    .B(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2834_ (.I(\minimax.regS_uc[12] ),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2835_ (.A1(_0278_),
    .A2(_0127_),
    .A3(_0275_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2836_ (.A1(_1856_),
    .A2(_1857_),
    .A3(_1858_),
    .A4(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2837_ (.A1(\minimax.regS_uc[12] ),
    .A2(_0219_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2838_ (.A1(_0187_),
    .A2(_0275_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2839_ (.A1(_1739_),
    .A2(_0276_),
    .B1(_0281_),
    .B2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2840_ (.A1(_0277_),
    .A2(_0280_),
    .A3(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2841_ (.A1(_0203_),
    .A2(_0273_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _2842_ (.A1(_0203_),
    .A2(_0273_),
    .A3(_0284_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2843_ (.A1(_0271_),
    .A2(net5),
    .B(_0285_),
    .C(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2844_ (.I(_0238_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2845_ (.A1(_0288_),
    .A2(net5),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2846_ (.I(_2017_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2847_ (.A1(_0277_),
    .A2(_0280_),
    .A3(_0283_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2848_ (.I(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2849_ (.A1(_2017_),
    .A2(_0272_),
    .A3(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2850_ (.A1(_0290_),
    .A2(_0292_),
    .B(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2851_ (.A1(_0203_),
    .A2(_0288_),
    .A3(net5),
    .A4(_0284_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2852_ (.A1(_0102_),
    .A2(_0218_),
    .A3(_0229_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2853_ (.I(_2049_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2854_ (.A1(_0238_),
    .A2(_0211_),
    .A3(_0272_),
    .A4(_0291_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2855_ (.A1(_0297_),
    .A2(_0242_),
    .A3(_0244_),
    .A4(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _2856_ (.A1(_0289_),
    .A2(_0294_),
    .B1(_0295_),
    .B2(_0296_),
    .C(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _2857_ (.A1(_0287_),
    .A2(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2858_ (.A1(_1876_),
    .A2(_1639_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2859_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2860_ (.A1(_0253_),
    .A2(_0270_),
    .B(_0301_),
    .C(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _2861_ (.A1(_0154_),
    .A2(_0252_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _2862_ (.A1(_0266_),
    .A2(_0269_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2863_ (.A1(_0287_),
    .A2(_0300_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2864_ (.A1(_0303_),
    .A2(_0305_),
    .A3(_0306_),
    .A4(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2865_ (.A1(_0231_),
    .A2(_0246_),
    .A3(_0250_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2866_ (.A1(_0102_),
    .A2(_0099_),
    .A3(_0218_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2867_ (.A1(_0162_),
    .A2(_0193_),
    .B(_0290_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2868_ (.A1(_0170_),
    .A2(_0090_),
    .A3(_0091_),
    .A4(_0196_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2869_ (.A1(_2071_),
    .A2(_0090_),
    .A3(_0091_),
    .A4(_0185_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2870_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0312_),
    .A4(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2871_ (.A1(_0310_),
    .A2(_0311_),
    .B(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2872_ (.I(_0196_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2873_ (.A1(_0193_),
    .A2(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2874_ (.A1(_0193_),
    .A2(_0316_),
    .B(_0170_),
    .C(_0161_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2875_ (.A1(_0297_),
    .A2(_0085_),
    .B1(_0317_),
    .B2(_0318_),
    .C(_0290_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2876_ (.A1(_0261_),
    .A2(_0315_),
    .A3(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2877_ (.A1(_0309_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2878_ (.A1(_0159_),
    .A2(_0183_),
    .B(_0309_),
    .C(_0320_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2879_ (.A1(_0254_),
    .A2(_0181_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2880_ (.I(_0259_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2881_ (.A1(_0254_),
    .A2(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2882_ (.I0(_0323_),
    .I1(_0325_),
    .S(_0177_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2883_ (.A1(_0231_),
    .A2(_0246_),
    .A3(_0250_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2884_ (.A1(_0261_),
    .A2(_0315_),
    .A3(_0319_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2885_ (.A1(_0326_),
    .A2(_0327_),
    .A3(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2886_ (.A1(_0154_),
    .A2(_0321_),
    .B(_0322_),
    .C(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2887_ (.A1(_2001_),
    .A2(_0152_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2888_ (.A1(_0159_),
    .A2(_0183_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2889_ (.A1(_0326_),
    .A2(_0327_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2890_ (.A1(_0254_),
    .A2(_0262_),
    .A3(_0309_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _2891_ (.A1(_0331_),
    .A2(_0332_),
    .A3(_0333_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2892_ (.A1(_0330_),
    .A2(_0335_),
    .B(_0302_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2893_ (.A1(_0304_),
    .A2(_0308_),
    .A3(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2894_ (.I(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2895_ (.A1(\bank1.rdata[0] ),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _2896_ (.A1(_0253_),
    .A2(_0270_),
    .B(_0307_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2897_ (.A1(_0305_),
    .A2(_0306_),
    .A3(_0301_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2898_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2899_ (.A1(_0330_),
    .A2(net373),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2900_ (.A1(_0340_),
    .A2(_0342_),
    .A3(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2901_ (.I(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2902_ (.A1(\bank3.rdata[0] ),
    .A2(_0345_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2903_ (.I(\bank2.rdata[0] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2904_ (.A1(net403),
    .A2(_0306_),
    .B(_0301_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2905_ (.A1(_0253_),
    .A2(_0270_),
    .A3(_0307_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2906_ (.A1(_0348_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2907_ (.I(_0350_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2908_ (.I(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2909_ (.A1(_0330_),
    .A2(net373),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2910_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2911_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2912_ (.I(_0340_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2913_ (.I(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2914_ (.I(_0341_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2915_ (.A1(\bank4.rdata[0] ),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2916_ (.A1(_0347_),
    .A2(_0352_),
    .B(_0355_),
    .C(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2917_ (.I(_0208_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2918_ (.I(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2919_ (.A1(_0346_),
    .A2(_0360_),
    .B(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2920_ (.A1(_0339_),
    .A2(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2921_ (.I(_0364_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2922_ (.I(\bank2.rdata[16] ),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2923_ (.I(_0350_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2924_ (.I(_0353_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2925_ (.I(_0356_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2926_ (.I(_0342_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2927_ (.A1(\bank4.rdata[16] ),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2928_ (.A1(_0365_),
    .A2(_0366_),
    .B(_0367_),
    .C(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2929_ (.A1(\bank3.rdata[16] ),
    .A2(_0345_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _2930_ (.I(_0361_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2931_ (.A1(_0371_),
    .A2(_0372_),
    .B(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2932_ (.I(_0337_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2933_ (.I(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2934_ (.A1(\bank1.rdata[16] ),
    .A2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2935_ (.A1(_0374_),
    .A2(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2936_ (.I(_0378_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2937_ (.I(\minimax.pc_fetch[1] ),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2938_ (.I0(net71),
    .I1(net78),
    .S(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2939_ (.I(_0380_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2940_ (.I(\bank2.rdata[1] ),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2941_ (.A1(\bank4.rdata[1] ),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2942_ (.A1(_0381_),
    .A2(_0352_),
    .B(_0355_),
    .C(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2943_ (.I(_0344_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2944_ (.A1(\bank3.rdata[1] ),
    .A2(_0384_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2945_ (.I(_0208_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2946_ (.A1(_0383_),
    .A2(_0385_),
    .B(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2947_ (.I(_0337_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2948_ (.A1(\bank1.rdata[1] ),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _2949_ (.A1(_0387_),
    .A2(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _2950_ (.I(_0390_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2951_ (.I(\bank2.rdata[17] ),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2952_ (.I(_0350_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2953_ (.I(_0353_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2954_ (.I(_0356_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2955_ (.I(_0342_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2956_ (.A1(\bank4.rdata[17] ),
    .A2(_0394_),
    .A3(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2957_ (.A1(_0391_),
    .A2(_0392_),
    .B(_0393_),
    .C(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2958_ (.I(_0344_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2959_ (.A1(\bank3.rdata[17] ),
    .A2(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2960_ (.A1(_0397_),
    .A2(_0399_),
    .B(_0362_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2961_ (.I(_0337_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2962_ (.A1(\bank1.rdata[17] ),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2963_ (.A1(_0400_),
    .A2(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2964_ (.I(_0403_),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2965_ (.I0(net82),
    .I1(net79),
    .S(_0379_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2966_ (.I(_0404_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2967_ (.I(\bank2.rdata[2] ),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2968_ (.A1(\bank4.rdata[2] ),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2969_ (.A1(_0405_),
    .A2(_0366_),
    .B(_0367_),
    .C(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2970_ (.A1(\bank3.rdata[2] ),
    .A2(_0345_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2971_ (.I(_0361_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2972_ (.A1(_0407_),
    .A2(_0408_),
    .B(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2973_ (.A1(\bank1.rdata[2] ),
    .A2(_0338_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2974_ (.A1(_0410_),
    .A2(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _2975_ (.I(_0412_),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2976_ (.I(\bank2.rdata[18] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2977_ (.A1(\bank4.rdata[18] ),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2978_ (.A1(_0413_),
    .A2(_0392_),
    .B(_0393_),
    .C(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2979_ (.A1(\bank3.rdata[18] ),
    .A2(_0384_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2980_ (.A1(_0415_),
    .A2(_0416_),
    .B(_0362_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2981_ (.A1(\bank1.rdata[18] ),
    .A2(_0401_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2982_ (.A1(_0417_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2983_ (.I(_0419_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2984_ (.I(\minimax.pc_fetch[1] ),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2985_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2986_ (.I0(net93),
    .I1(net80),
    .S(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2987_ (.I(_0422_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2988_ (.I(\bank2.rdata[3] ),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _2989_ (.I(_0350_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2990_ (.I(_0353_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2991_ (.A1(\bank4.rdata[3] ),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2992_ (.A1(_0423_),
    .A2(_0424_),
    .B(_0425_),
    .C(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2993_ (.I(_0344_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2994_ (.A1(\bank3.rdata[3] ),
    .A2(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2995_ (.A1(_0427_),
    .A2(_0429_),
    .B(_0373_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2996_ (.I(_0375_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2997_ (.A1(\bank1.rdata[3] ),
    .A2(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2998_ (.A1(_0430_),
    .A2(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _2999_ (.I(_0433_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3000_ (.I(\bank1.rdata[19] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3001_ (.A1(_0352_),
    .A2(_0355_),
    .B(_0303_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3002_ (.I(_0353_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3003_ (.A1(_0348_),
    .A2(net396),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3004_ (.I0(\bank3.rdata[19] ),
    .I1(\bank4.rdata[19] ),
    .S(_0436_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3005_ (.A1(_0340_),
    .A2(_0341_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3006_ (.I(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3007_ (.A1(\bank2.rdata[19] ),
    .A2(_0437_),
    .B1(_0438_),
    .B2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3008_ (.I(_0303_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3009_ (.A1(_0434_),
    .A2(_0435_),
    .B1(_0441_),
    .B2(_0442_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3010_ (.I0(net96),
    .I1(net81),
    .S(_0421_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3011_ (.I(_0443_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3012_ (.I(\bank2.rdata[4] ),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3013_ (.A1(\bank4.rdata[4] ),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3014_ (.A1(_0444_),
    .A2(_0424_),
    .B(_0367_),
    .C(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3015_ (.A1(\bank3.rdata[4] ),
    .A2(_0345_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3016_ (.A1(_0446_),
    .A2(_0447_),
    .B(_0373_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3017_ (.A1(\bank1.rdata[4] ),
    .A2(_0431_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3018_ (.A1(_0448_),
    .A2(_0449_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3019_ (.I(_0450_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3020_ (.I(\bank2.rdata[20] ),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3021_ (.A1(\bank4.rdata[20] ),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3022_ (.A1(_0451_),
    .A2(_0392_),
    .B(_0355_),
    .C(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3023_ (.A1(\bank3.rdata[20] ),
    .A2(_0384_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3024_ (.A1(_0453_),
    .A2(_0454_),
    .B(_0362_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3025_ (.A1(\bank1.rdata[20] ),
    .A2(_0401_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3026_ (.A1(_0455_),
    .A2(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3027_ (.I(_0457_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3028_ (.I0(net97),
    .I1(net83),
    .S(_0421_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3029_ (.I(_0458_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3030_ (.I(\bank2.rdata[5] ),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3031_ (.I(_0350_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3032_ (.I(_0356_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3033_ (.I(_0342_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3034_ (.A1(\bank4.rdata[5] ),
    .A2(_0461_),
    .A3(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3035_ (.A1(_0459_),
    .A2(_0460_),
    .B(_0425_),
    .C(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3036_ (.A1(\bank3.rdata[5] ),
    .A2(_0428_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3037_ (.A1(_0464_),
    .A2(_0465_),
    .B(_0209_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3038_ (.A1(\bank1.rdata[5] ),
    .A2(_0431_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3039_ (.A1(_0466_),
    .A2(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3040_ (.I(_0468_),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3041_ (.I(\bank2.rdata[21] ),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3042_ (.A1(\bank4.rdata[21] ),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3043_ (.A1(_0469_),
    .A2(_0352_),
    .B(_0355_),
    .C(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3044_ (.A1(\bank3.rdata[21] ),
    .A2(_0384_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3045_ (.A1(_0471_),
    .A2(_0472_),
    .B(_0386_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3046_ (.A1(\bank1.rdata[21] ),
    .A2(_0388_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _3047_ (.A1(_0473_),
    .A2(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _3048_ (.I(_0475_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3049_ (.I0(net98),
    .I1(net84),
    .S(_0421_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3050_ (.I(_0476_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3051_ (.I(\bank2.rdata[6] ),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3052_ (.A1(\bank4.rdata[6] ),
    .A2(_0461_),
    .A3(_0462_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3053_ (.A1(_0477_),
    .A2(_0424_),
    .B(_0425_),
    .C(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3054_ (.A1(\bank3.rdata[6] ),
    .A2(_0428_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3055_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0209_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3056_ (.A1(\bank1.rdata[6] ),
    .A2(_0431_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3057_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3058_ (.I(_0483_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3059_ (.I(\bank1.rdata[22] ),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3060_ (.I0(\bank3.rdata[22] ),
    .I1(\bank4.rdata[22] ),
    .S(_0436_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3061_ (.A1(\bank2.rdata[22] ),
    .A2(_0437_),
    .B1(_0485_),
    .B2(_0440_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3062_ (.A1(_0484_),
    .A2(_0435_),
    .B1(_0486_),
    .B2(_0442_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3063_ (.I0(net99),
    .I1(net85),
    .S(_0421_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3064_ (.I(_0487_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3065_ (.I(\bank2.rdata[7] ),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3066_ (.A1(\bank4.rdata[7] ),
    .A2(_0461_),
    .A3(_0462_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3067_ (.A1(_0488_),
    .A2(_0424_),
    .B(_0425_),
    .C(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3068_ (.A1(\bank3.rdata[7] ),
    .A2(_0428_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3069_ (.A1(_0490_),
    .A2(_0491_),
    .B(_0209_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3070_ (.A1(\bank1.rdata[7] ),
    .A2(_0376_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3071_ (.A1(_0492_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3072_ (.I(_0494_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3073_ (.I(\bank2.rdata[23] ),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3074_ (.A1(\bank4.rdata[23] ),
    .A2(_0356_),
    .A3(_0342_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3075_ (.A1(_0495_),
    .A2(_0352_),
    .B(_0436_),
    .C(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3076_ (.A1(\bank3.rdata[23] ),
    .A2(_0384_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3077_ (.A1(_0497_),
    .A2(_0498_),
    .B(_0386_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3078_ (.A1(\bank1.rdata[23] ),
    .A2(_0375_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3079_ (.A1(_0499_),
    .A2(_0500_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3080_ (.I(_0501_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3081_ (.I(_0420_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3082_ (.I0(net100),
    .I1(net86),
    .S(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3083_ (.I(_0503_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3084_ (.I(\bank2.rdata[8] ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3085_ (.I(_0354_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3086_ (.A1(\bank4.rdata[8] ),
    .A2(_0461_),
    .A3(_0462_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3087_ (.A1(_0504_),
    .A2(_0460_),
    .B(_0505_),
    .C(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3088_ (.I(_0344_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3089_ (.A1(\bank3.rdata[8] ),
    .A2(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3090_ (.A1(_0507_),
    .A2(_0509_),
    .B(_0209_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3091_ (.I(_0337_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3092_ (.A1(\bank1.rdata[8] ),
    .A2(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _3093_ (.A1(_0510_),
    .A2(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3094_ (.I(_0513_),
    .ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3095_ (.A1(_0361_),
    .A2(_0343_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3096_ (.A1(\bank4.rdata[24] ),
    .A2(_0348_),
    .A3(_0349_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3097_ (.A1(\bank2.rdata[24] ),
    .A2(_0460_),
    .B(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3098_ (.A1(_0304_),
    .A2(_0308_),
    .B(\bank3.rdata[24] ),
    .C(_0505_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3099_ (.A1(\bank1.rdata[24] ),
    .A2(_0401_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3100_ (.A1(_0514_),
    .A2(_0516_),
    .B(_0517_),
    .C(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3101_ (.I(_0519_),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3102_ (.A1(_0379_),
    .A2(net87),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3103_ (.A1(_0379_),
    .A2(_0513_),
    .B(_0520_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3104_ (.I(\bank2.rdata[9] ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3105_ (.A1(\bank4.rdata[9] ),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3106_ (.A1(_0521_),
    .A2(_0366_),
    .B(_0367_),
    .C(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3107_ (.A1(\bank3.rdata[9] ),
    .A2(_0345_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3108_ (.A1(_0523_),
    .A2(_0524_),
    .B(_0373_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3109_ (.A1(\bank1.rdata[9] ),
    .A2(_0376_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3110_ (.A1(_0525_),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3111_ (.I(_0527_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3112_ (.I(\bank1.rdata[25] ),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3113_ (.I0(\bank3.rdata[25] ),
    .I1(\bank4.rdata[25] ),
    .S(_0354_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3114_ (.A1(\bank2.rdata[25] ),
    .A2(_0437_),
    .B1(_0529_),
    .B2(_0440_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3115_ (.A1(_0528_),
    .A2(_0435_),
    .B1(_0530_),
    .B2(_0442_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3116_ (.I0(net102),
    .I1(net88),
    .S(_0502_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3117_ (.I(_0531_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3118_ (.I(\bank2.rdata[10] ),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3119_ (.A1(\bank4.rdata[10] ),
    .A2(_0394_),
    .A3(_0395_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3120_ (.A1(_0532_),
    .A2(_0366_),
    .B(_0367_),
    .C(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3121_ (.A1(\bank3.rdata[10] ),
    .A2(_0398_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3122_ (.A1(_0534_),
    .A2(_0535_),
    .B(_0409_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3123_ (.A1(\bank1.rdata[10] ),
    .A2(_0338_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3124_ (.A1(_0536_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3125_ (.I(_0538_),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3126_ (.A1(\bank1.rdata[26] ),
    .A2(_0388_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3127_ (.I0(\bank2.rdata[26] ),
    .I1(\bank4.rdata[26] ),
    .S(_0351_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3128_ (.A1(\bank3.rdata[26] ),
    .A2(_0386_),
    .A3(_0508_),
    .B1(_0540_),
    .B2(net402),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3129_ (.A1(_0539_),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3130_ (.I(_0542_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3131_ (.I0(net72),
    .I1(net89),
    .S(_0502_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3132_ (.I(_0543_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3133_ (.I(\bank2.rdata[11] ),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3134_ (.A1(\bank4.rdata[11] ),
    .A2(_0394_),
    .A3(_0395_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3135_ (.A1(_0544_),
    .A2(_0366_),
    .B(_0393_),
    .C(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3136_ (.A1(\bank3.rdata[11] ),
    .A2(_0398_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3137_ (.A1(_0546_),
    .A2(_0547_),
    .B(_0409_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3138_ (.A1(\bank1.rdata[11] ),
    .A2(_0338_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3139_ (.A1(_0548_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3140_ (.I(_0550_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3141_ (.I(\bank1.rdata[27] ),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3142_ (.I0(\bank3.rdata[27] ),
    .I1(\bank4.rdata[27] ),
    .S(_0436_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3143_ (.A1(\bank2.rdata[27] ),
    .A2(_0437_),
    .B1(_0552_),
    .B2(_0440_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3144_ (.A1(_0551_),
    .A2(_0435_),
    .B1(_0553_),
    .B2(_0442_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3145_ (.I0(net73),
    .I1(net90),
    .S(_0502_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3146_ (.I(_0554_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3147_ (.I(\bank2.rdata[12] ),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3148_ (.A1(\bank4.rdata[12] ),
    .A2(_0394_),
    .A3(_0395_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3149_ (.A1(_0555_),
    .A2(_0392_),
    .B(_0393_),
    .C(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3150_ (.A1(\bank3.rdata[12] ),
    .A2(_0398_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3151_ (.A1(_0557_),
    .A2(_0558_),
    .B(_0409_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3152_ (.A1(\bank1.rdata[12] ),
    .A2(_0338_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3153_ (.A1(_0559_),
    .A2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3154_ (.I(_0561_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3155_ (.A1(\bank1.rdata[28] ),
    .A2(_0388_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3156_ (.I0(\bank2.rdata[28] ),
    .I1(\bank4.rdata[28] ),
    .S(_0351_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3157_ (.A1(\bank3.rdata[28] ),
    .A2(_0361_),
    .A3(_0508_),
    .B1(_0563_),
    .B2(net402),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _3158_ (.A1(_0562_),
    .A2(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3159_ (.I(_0565_),
    .ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3160_ (.I0(net74),
    .I1(net91),
    .S(_0502_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3161_ (.I(_0566_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3162_ (.I(\bank2.rdata[13] ),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3163_ (.A1(\bank4.rdata[13] ),
    .A2(_0394_),
    .A3(_0395_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3164_ (.A1(_0567_),
    .A2(_0392_),
    .B(_0393_),
    .C(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3165_ (.A1(\bank3.rdata[13] ),
    .A2(_0398_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3166_ (.A1(_0569_),
    .A2(_0570_),
    .B(_0409_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3167_ (.A1(\bank1.rdata[13] ),
    .A2(_0401_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3168_ (.A1(_0571_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3169_ (.I(_0573_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3170_ (.A1(\bank4.rdata[29] ),
    .A2(_0348_),
    .A3(_0349_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3171_ (.A1(\bank2.rdata[29] ),
    .A2(_0460_),
    .B(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3172_ (.A1(\bank3.rdata[29] ),
    .A2(_0386_),
    .A3(_0508_),
    .B1(_0388_),
    .B2(\bank1.rdata[29] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3173_ (.A1(_0514_),
    .A2(_0575_),
    .B(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3174_ (.I(_0577_),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3175_ (.I0(net75),
    .I1(net92),
    .S(_0420_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3176_ (.I(_0578_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3177_ (.I(\bank2.rdata[14] ),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3178_ (.A1(\bank4.rdata[14] ),
    .A2(_0461_),
    .A3(_0462_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3179_ (.A1(_0579_),
    .A2(_0424_),
    .B(_0425_),
    .C(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3180_ (.A1(\bank3.rdata[14] ),
    .A2(_0428_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3181_ (.A1(_0581_),
    .A2(_0582_),
    .B(_0373_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3182_ (.A1(\bank1.rdata[14] ),
    .A2(_0376_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3183_ (.A1(_0583_),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3184_ (.I(_0585_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3185_ (.I(\bank1.rdata[30] ),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3186_ (.I0(\bank3.rdata[30] ),
    .I1(\bank4.rdata[30] ),
    .S(_0354_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3187_ (.A1(\bank2.rdata[30] ),
    .A2(_0437_),
    .B1(_0587_),
    .B2(_0440_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3188_ (.A1(_0586_),
    .A2(_0435_),
    .B1(_0588_),
    .B2(_0442_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3189_ (.I0(net76),
    .I1(net94),
    .S(_0420_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3190_ (.I(_0589_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3191_ (.I0(\bank2.rdata[15] ),
    .I1(\bank4.rdata[15] ),
    .S(_0351_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3192_ (.A1(\bank3.rdata[15] ),
    .A2(_0362_),
    .A3(_0508_),
    .B1(_0590_),
    .B2(net402),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3193_ (.A1(\bank1.rdata[15] ),
    .A2(_0376_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3194_ (.A1(_0591_),
    .A2(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3195_ (.I(_0593_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3196_ (.A1(_0439_),
    .A2(_0514_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3197_ (.I0(\bank3.rdata[31] ),
    .I1(\bank4.rdata[31] ),
    .S(_0354_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3198_ (.A1(_0303_),
    .A2(_0351_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3199_ (.A1(\bank2.rdata[31] ),
    .A2(_0594_),
    .B1(_0595_),
    .B2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3200_ (.A1(\bank1.rdata[31] ),
    .A2(_0375_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _3201_ (.A1(_0597_),
    .A2(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3202_ (.I(_0599_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3203_ (.I0(net77),
    .I1(net95),
    .S(_0420_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3204_ (.I(_0600_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3205_ (.I0(\minimax.regD_ex[4] ),
    .I1(\minimax.regD_uc[4] ),
    .S(_1733_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3206_ (.I(_0601_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _3207_ (.I0(\minimax.regD_ex[5] ),
    .I1(\minimax.regD_uc[5] ),
    .S(_1733_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3208_ (.I(_0602_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _3209_ (.I0(\minimax.regD_ex[6] ),
    .I1(\minimax.regD_uc[6] ),
    .S(_2034_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3210_ (.I(_0603_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3211_ (.I0(\minimax.regD_ex[13] ),
    .I1(\minimax.regD_uc[13] ),
    .S(_1730_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3212_ (.I(_0604_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3213_ (.I0(\minimax.regD_ex[14] ),
    .I1(\minimax.regD_uc[14] ),
    .S(_1728_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3214_ (.I(_0605_),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3215_ (.A1(\minimax.regD_uc[15] ),
    .A2(_1856_),
    .A3(_1857_),
    .A4(_1858_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3216_ (.A1(\minimax.regD_ex[15] ),
    .A2(_1868_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3217_ (.A1(_1856_),
    .A2(_1858_),
    .B(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3218_ (.A1(\minimax.regD_uc[15] ),
    .A2(_1737_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3219_ (.A1(_1857_),
    .A2(_0607_),
    .B(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3220_ (.A1(_0606_),
    .A2(_0608_),
    .A3(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3221_ (.I(_0611_),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3222_ (.I0(\minimax.regD_ex[16] ),
    .I1(\minimax.regD_uc[16] ),
    .S(_1729_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3223_ (.I(_0612_),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3224_ (.I(_1729_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3225_ (.I0(\minimax.regD_ex[17] ),
    .I1(\minimax.regD_uc[17] ),
    .S(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3226_ (.I(_0614_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3227_ (.I0(\minimax.regD_ex[18] ),
    .I1(\minimax.regD_uc[18] ),
    .S(_1730_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3228_ (.I(_0615_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3229_ (.I0(\minimax.regD_ex[19] ),
    .I1(\minimax.regD_uc[19] ),
    .S(_0613_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3230_ (.I(_0616_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3231_ (.I0(\minimax.regD_ex[20] ),
    .I1(\minimax.regD_uc[20] ),
    .S(_0613_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3232_ (.I(_0617_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3233_ (.I0(\minimax.regD_ex[21] ),
    .I1(\minimax.regD_uc[21] ),
    .S(_1729_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3234_ (.I(_0618_),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3235_ (.I0(\minimax.regD_ex[22] ),
    .I1(\minimax.regD_uc[22] ),
    .S(_1730_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3236_ (.I(_0619_),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3237_ (.I0(\minimax.regD_ex[23] ),
    .I1(\minimax.regD_uc[23] ),
    .S(_0613_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3238_ (.I(_0620_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3239_ (.I0(\minimax.regD_ex[24] ),
    .I1(\minimax.regD_uc[24] ),
    .S(_0613_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3240_ (.I(_0621_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3241_ (.I0(\minimax.regD_ex[25] ),
    .I1(\minimax.regD_uc[25] ),
    .S(_1730_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3242_ (.I(_0622_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3243_ (.I0(\minimax.regD_ex[26] ),
    .I1(\minimax.regD_uc[26] ),
    .S(_1731_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3244_ (.I(_0623_),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3245_ (.I0(\minimax.regD_ex[27] ),
    .I1(\minimax.regD_uc[27] ),
    .S(_1731_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3246_ (.I(_0624_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3247_ (.I0(\minimax.regD_ex[28] ),
    .I1(\minimax.regD_uc[28] ),
    .S(_1732_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _3248_ (.I(_0625_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3249_ (.I0(\minimax.regD_ex[29] ),
    .I1(\minimax.regD_uc[29] ),
    .S(_1731_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3250_ (.I(_0626_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3251_ (.I0(\minimax.regD_ex[30] ),
    .I1(\minimax.regD_uc[30] ),
    .S(_1732_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3252_ (.I(_0627_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3253_ (.I0(\minimax.regD_ex[31] ),
    .I1(\minimax.regD_uc[31] ),
    .S(_1731_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3254_ (.I(_0628_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3256_ (.A1(\bank4.was_en ),
    .A2(_0596_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3257_ (.A1(_0505_),
    .A2(_0629_),
    .B(net363),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3258_ (.I(_0630_),
    .Z(\bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3259_ (.A1(\bank3.was_en ),
    .A2(_0505_),
    .A3(_0596_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3260_ (.A1(net362),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3261_ (.I(_0632_),
    .Z(\bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3262_ (.A1(\bank2.was_en ),
    .A2(_0594_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3263_ (.A1(net361),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3264_ (.I(_0634_),
    .Z(\bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3265_ (.A1(net399),
    .A2(net392),
    .A3(_1692_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3266_ (.A1(_1632_),
    .A2(_0635_),
    .ZN(\bank1.wen_mask[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3267_ (.A1(\bank1.was_en ),
    .A2(_0431_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3268_ (.A1(net360),
    .A2(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3269_ (.I(_0637_),
    .Z(\bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3270_ (.I(_0290_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3271_ (.I(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3272_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3273_ (.I(net376),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3274_ (.A1(_1654_),
    .A2(_1759_),
    .B(_1649_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3275_ (.I0(_0641_),
    .I1(_0642_),
    .S(_1849_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3276_ (.A1(_1851_),
    .A2(_1638_),
    .A3(_1696_),
    .A4(_1660_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3277_ (.A1(_1812_),
    .A2(_1847_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3278_ (.A1(_0643_),
    .A2(_0644_),
    .B1(_0645_),
    .B2(net394),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3279_ (.A1(_1809_),
    .A2(_0640_),
    .A3(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3280_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3281_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3282_ (.A1(_1735_),
    .A2(_1823_),
    .B(_1832_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3283_ (.I(_0165_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3284_ (.A1(_0651_),
    .A2(_1870_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3285_ (.A1(_1846_),
    .A2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3286_ (.I(_0190_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3287_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3288_ (.I(_0655_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3289_ (.I(_0191_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3290_ (.A1(_0656_),
    .A2(_1859_),
    .B1(_1853_),
    .B2(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3291_ (.A1(_0650_),
    .A2(_0653_),
    .A3(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3292_ (.A1(\minimax.dly16_lwsp ),
    .A2(\minimax.dly16_lw ),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _3293_ (.I(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3294_ (.I(_0234_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3295_ (.A1(_0662_),
    .A2(_1763_),
    .A3(_0641_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3296_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3297_ (.A1(_1774_),
    .A2(_0645_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3298_ (.A1(_1655_),
    .A2(_0635_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3299_ (.A1(_1650_),
    .A2(_1779_),
    .A3(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3300_ (.A1(_2043_),
    .A2(_1654_),
    .A3(net397),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3301_ (.A1(_1849_),
    .A2(_0665_),
    .B1(_0667_),
    .B2(_0668_),
    .C(_0657_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3302_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3303_ (.A1(_1638_),
    .A2(_1660_),
    .A3(_0635_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3304_ (.A1(_1716_),
    .A2(_1720_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3305_ (.A1(_1650_),
    .A2(_0671_),
    .A3(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3306_ (.I(_0232_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3307_ (.A1(_0674_),
    .A2(_1939_),
    .A3(_0235_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3308_ (.A1(_0673_),
    .A2(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3309_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3310_ (.I(_0232_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3311_ (.A1(_0678_),
    .A2(_0233_),
    .A3(_0235_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3312_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3313_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3314_ (.A1(_0234_),
    .A2(_1771_),
    .A3(_1674_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3315_ (.I(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3316_ (.A1(_0650_),
    .A2(_0658_),
    .A3(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3317_ (.A1(_0650_),
    .A2(_0681_),
    .B(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3318_ (.A1(_0674_),
    .A2(_1939_),
    .A3(_0109_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3319_ (.A1(_1779_),
    .A2(_0666_),
    .B(_0671_),
    .C(_1649_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3320_ (.A1(_0675_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3321_ (.A1(_0686_),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3322_ (.A1(_0650_),
    .A2(_0689_),
    .B(_0658_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3323_ (.A1(_0677_),
    .A2(_0685_),
    .B(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3324_ (.A1(_1881_),
    .A2(_0664_),
    .B1(_0670_),
    .B2(\minimax.pc_fetch_dly[1] ),
    .C(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3325_ (.A1(_0649_),
    .A2(_0659_),
    .B1(_0661_),
    .B2(_0390_),
    .C(_0692_),
    .ZN(\minimax.aluX[1] ));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _3326_ (.A1(_1809_),
    .A2(_0639_),
    .A3(_0646_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3327_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3328_ (.I(_0694_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3329_ (.I(_0686_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3330_ (.I(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3331_ (.I(_1811_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3332_ (.I(_0179_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3333_ (.A1(\minimax.regS_ex[2] ),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3334_ (.A1(_1777_),
    .A2(_0699_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3335_ (.A1(_0698_),
    .A2(_1757_),
    .B(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3336_ (.I(_0682_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(_1881_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3338_ (.A1(_0702_),
    .A2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3339_ (.A1(_0697_),
    .A2(_0702_),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3340_ (.A1(_0675_),
    .A2(_0679_),
    .A3(_0687_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3341_ (.A1(_0707_),
    .A2(_0702_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3342_ (.A1(_0673_),
    .A2(_0675_),
    .A3(_0706_),
    .B1(_0708_),
    .B2(_1881_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3343_ (.I(_0663_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3344_ (.I(_0669_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3345_ (.A1(_1895_),
    .A2(_0710_),
    .B1(_0711_),
    .B2(\minimax.pc_fetch_dly[2] ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(_0709_),
    .A2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3347_ (.A1(_1874_),
    .A2(_0695_),
    .B(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3348_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0661_),
    .B(_0714_),
    .ZN(\minimax.aluX[2] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3349_ (.A1(\minimax.dly16_lwsp ),
    .A2(\minimax.dly16_lw ),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3350_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3351_ (.A1(\bank1.rdata[3] ),
    .A2(_0511_),
    .B(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3352_ (.I(_0663_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3353_ (.I(_0676_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3354_ (.I(_0288_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3355_ (.I(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3356_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3357_ (.A1(_0195_),
    .A2(_1889_),
    .B(_1893_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3358_ (.A1(_0722_),
    .A2(_1890_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3359_ (.A1(_0234_),
    .A2(_1674_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3360_ (.A1(_1763_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3361_ (.A1(_1902_),
    .A2(_0696_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3362_ (.A1(_0724_),
    .A2(_1902_),
    .A3(_0726_),
    .B(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3363_ (.A1(_0719_),
    .A2(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3364_ (.I(_0707_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3365_ (.A1(_1902_),
    .A2(_0730_),
    .B(_0724_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3366_ (.A1(_1977_),
    .A2(_0718_),
    .B1(_0729_),
    .B2(_0731_),
    .C1(_0711_),
    .C2(\minimax.pc_fetch_dly[3] ),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3367_ (.A1(_1912_),
    .A2(_0649_),
    .B1(_0717_),
    .B2(_0430_),
    .C(_0732_),
    .ZN(\minimax.aluX[3] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3368_ (.A1(\bank1.rdata[4] ),
    .A2(_0511_),
    .B(_0716_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3369_ (.A1(_2007_),
    .A2(_0696_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3370_ (.A1(_1976_),
    .A2(_2007_),
    .A3(_0726_),
    .B(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3371_ (.A1(_0719_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3372_ (.A1(_2007_),
    .A2(_0730_),
    .B(_1976_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3373_ (.A1(_1966_),
    .A2(_0718_),
    .B1(_0736_),
    .B2(_0737_),
    .C1(_0711_),
    .C2(\minimax.pc_fetch_dly[4] ),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3374_ (.A1(_1959_),
    .A2(_0649_),
    .B1(_0733_),
    .B2(_0448_),
    .C(_0738_),
    .ZN(\minimax.aluX[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3375_ (.I(_0375_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3376_ (.I(_0715_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3377_ (.I(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3378_ (.A1(\bank1.rdata[5] ),
    .A2(_0739_),
    .B(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3379_ (.I(_0726_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3380_ (.I(_0686_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3381_ (.A1(_1994_),
    .A2(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3382_ (.A1(_1965_),
    .A2(_1994_),
    .A3(_0743_),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3383_ (.A1(_0677_),
    .A2(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3384_ (.A1(_1994_),
    .A2(_0730_),
    .B(_1965_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3385_ (.A1(_2037_),
    .A2(_0718_),
    .B1(_0747_),
    .B2(_0748_),
    .C1(_0711_),
    .C2(\minimax.pc_fetch_dly[5] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3386_ (.A1(_1981_),
    .A2(_0695_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3387_ (.A1(_0466_),
    .A2(_0742_),
    .B(_0749_),
    .C(_0750_),
    .ZN(\minimax.aluX[5] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3388_ (.A1(\bank1.rdata[6] ),
    .A2(_0739_),
    .B(_0741_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3389_ (.A1(_2037_),
    .A2(_2015_),
    .A3(_0703_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3390_ (.A1(_2015_),
    .A2(_0681_),
    .B(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3391_ (.I(_0689_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3392_ (.A1(_2015_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3393_ (.A1(_0677_),
    .A2(_0753_),
    .B1(_0755_),
    .B2(_2006_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3394_ (.A1(_0115_),
    .A2(_0664_),
    .B1(_0670_),
    .B2(\minimax.pc_fetch_dly[6] ),
    .C(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3395_ (.I(_0693_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3396_ (.A1(_2031_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3397_ (.A1(_0481_),
    .A2(_0751_),
    .B(_0757_),
    .C(_0759_),
    .ZN(\minimax.aluX[6] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3398_ (.A1(\bank1.rdata[7] ),
    .A2(_0739_),
    .B(_0741_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3399_ (.A1(_0146_),
    .A2(_0703_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3400_ (.A1(_0146_),
    .A2(_0680_),
    .B1(_0761_),
    .B2(_2047_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3401_ (.A1(_0146_),
    .A2(_0689_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3402_ (.A1(_0719_),
    .A2(_0762_),
    .B1(_0763_),
    .B2(_2047_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3403_ (.A1(_0170_),
    .A2(_0664_),
    .B1(_0670_),
    .B2(\minimax.pc_fetch_dly[7] ),
    .C(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3404_ (.A1(_2064_),
    .A2(_0758_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3405_ (.A1(_0492_),
    .A2(_0760_),
    .B(_0765_),
    .C(_0766_),
    .ZN(\minimax.aluX[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3406_ (.I(_0660_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3407_ (.A1(_0170_),
    .A2(_0162_),
    .A3(_0703_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3408_ (.A1(_0162_),
    .A2(_0681_),
    .B(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3409_ (.A1(_0162_),
    .A2(_0689_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3410_ (.A1(_0719_),
    .A2(_0769_),
    .B1(_0770_),
    .B2(_0107_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3411_ (.A1(_0316_),
    .A2(_0664_),
    .B1(_0670_),
    .B2(\minimax.pc_fetch_dly[8] ),
    .C(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3412_ (.A1(_0119_),
    .A2(_0758_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3413_ (.A1(_0513_),
    .A2(_0767_),
    .B(_0772_),
    .C(_0773_),
    .ZN(\minimax.aluX[8] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3414_ (.A1(\bank1.rdata[9] ),
    .A2(_0511_),
    .B(_0716_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(_0316_),
    .A2(_0754_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3416_ (.A1(_0316_),
    .A2(_0680_),
    .B1(_0726_),
    .B2(_0317_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3417_ (.I(_0676_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3418_ (.A1(_0185_),
    .A2(_0775_),
    .B1(_0776_),
    .B2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3419_ (.A1(net3),
    .A2(_0718_),
    .B1(_0711_),
    .B2(\minimax.pc_fetch_dly[9] ),
    .C(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3420_ (.A1(_0172_),
    .A2(_0649_),
    .B1(_0774_),
    .B2(_0525_),
    .C(_0779_),
    .ZN(\minimax.aluX[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3421_ (.I(_0710_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3422_ (.I(_0777_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3423_ (.I(_0726_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3424_ (.A1(_1871_),
    .A2(_0647_),
    .A3(_0697_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3425_ (.A1(_1871_),
    .A2(_1870_),
    .A3(_0782_),
    .B(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3426_ (.A1(_0781_),
    .A2(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3427_ (.A1(_0694_),
    .A2(_0754_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3428_ (.A1(_1871_),
    .A2(_0786_),
    .B(_1870_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3429_ (.A1(net13),
    .A2(_0780_),
    .B1(_0785_),
    .B2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3430_ (.A1(_0339_),
    .A2(_0363_),
    .A3(_0661_),
    .B(_0788_),
    .ZN(\minimax.aluX[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3431_ (.A1(_0207_),
    .A2(_0648_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3432_ (.I(_0680_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3433_ (.A1(_0720_),
    .A2(net3),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3434_ (.I(_0682_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3435_ (.A1(_0791_),
    .A2(_0324_),
    .A3(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3436_ (.A1(_0324_),
    .A2(_0790_),
    .B(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3437_ (.A1(_0324_),
    .A2(_0754_),
    .B(_0791_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3438_ (.A1(_0781_),
    .A2(_0794_),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3439_ (.A1(net4),
    .A2(_0780_),
    .B(_0789_),
    .C(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3440_ (.A1(_0536_),
    .A2(_0537_),
    .A3(_0661_),
    .B(_0797_),
    .ZN(\minimax.aluX[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3441_ (.I(_0660_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3442_ (.I(_0663_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3443_ (.I(_0693_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3444_ (.I(_0777_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3445_ (.A1(_0267_),
    .A2(_0217_),
    .A3(_0792_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3446_ (.A1(_0217_),
    .A2(_0681_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3447_ (.A1(_0217_),
    .A2(_0754_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3448_ (.A1(_0801_),
    .A2(_0803_),
    .B1(_0804_),
    .B2(_0213_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3449_ (.A1(net5),
    .A2(_0799_),
    .B1(_0800_),
    .B2(_0505_),
    .C(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3450_ (.A1(_0548_),
    .A2(_0549_),
    .A3(_0798_),
    .B(_0806_),
    .ZN(\minimax.aluX[11] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3451_ (.A1(_0292_),
    .A2(_0697_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3452_ (.A1(_0289_),
    .A2(_0292_),
    .A3(_0743_),
    .B(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3453_ (.A1(_0801_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3454_ (.A1(_0292_),
    .A2(_0730_),
    .B(_0289_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _3455_ (.A1(net6),
    .A2(_0799_),
    .B1(_0809_),
    .B2(_0810_),
    .C1(_0800_),
    .C2(_0460_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3456_ (.A1(_0559_),
    .A2(_0560_),
    .A3(_0798_),
    .B(_0811_),
    .ZN(\minimax.aluX[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3457_ (.I(_0647_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3458_ (.A1(_0315_),
    .A2(_0319_),
    .B(_0326_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3459_ (.A1(_0267_),
    .A2(_0268_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3460_ (.A1(_0267_),
    .A2(_0248_),
    .A3(_0249_),
    .A4(_0237_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3461_ (.A1(_0815_),
    .A2(_0300_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3462_ (.A1(_0267_),
    .A2(_0268_),
    .B(_0261_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3463_ (.A1(_0813_),
    .A2(_0814_),
    .B(_0816_),
    .C(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3464_ (.A1(_0154_),
    .A2(_0252_),
    .B(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3465_ (.A1(_0287_),
    .A2(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3466_ (.I(_0271_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3467_ (.A1(_0821_),
    .A2(net6),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3468_ (.I(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3469_ (.I(_0203_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3470_ (.A1(_0075_),
    .A2(_2053_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3471_ (.I(_0257_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3472_ (.I0(\minimax.regS_ex[13] ),
    .I1(\minimax.regS_uc[13] ),
    .S(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3473_ (.A1(_1642_),
    .A2(_0825_),
    .B(_0827_),
    .C(_0128_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3474_ (.A1(_0240_),
    .A2(_0284_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3475_ (.A1(_0296_),
    .A2(_0829_),
    .B(_0828_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3476_ (.I(_0101_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3477_ (.A1(_1759_),
    .A2(_0825_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3478_ (.A1(\minimax.regS_ex[12] ),
    .A2(\minimax.regS_ex[13] ),
    .A3(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3479_ (.A1(\minimax.regS_uc[12] ),
    .A2(\minimax.regS_uc[13] ),
    .A3(_0832_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3480_ (.I0(_0833_),
    .I1(_0834_),
    .S(_0084_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3481_ (.A1(_0188_),
    .A2(_0272_),
    .A3(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3482_ (.A1(_2050_),
    .A2(_0242_),
    .A3(_0244_),
    .A4(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3483_ (.A1(_0831_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _3484_ (.A1(_0824_),
    .A2(_0828_),
    .B1(_0830_),
    .B2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3485_ (.A1(_0820_),
    .A2(_0823_),
    .A3(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3486_ (.A1(_0812_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3487_ (.A1(_0823_),
    .A2(_0828_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3488_ (.I0(_0744_),
    .I1(_0683_),
    .S(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3489_ (.I(_0777_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3490_ (.A1(_0823_),
    .A2(_0828_),
    .B1(_0843_),
    .B2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3491_ (.A1(net7),
    .A2(_0780_),
    .B(_0841_),
    .C(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3492_ (.A1(_0571_),
    .A2(_0572_),
    .A3(_0798_),
    .B(_0846_),
    .ZN(\minimax.aluX[13] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3493_ (.A1(\bank1.rdata[14] ),
    .A2(_0739_),
    .B(_0716_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3494_ (.A1(_0822_),
    .A2(_0839_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3495_ (.A1(net403),
    .A2(_0306_),
    .B(_0287_),
    .C(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3496_ (.A1(_0823_),
    .A2(_0839_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3497_ (.A1(_0300_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3498_ (.A1(_0823_),
    .A2(_0839_),
    .B(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3499_ (.A1(_0849_),
    .A2(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_0288_),
    .A2(net7),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3501_ (.A1(\minimax.regS_ex[14] ),
    .A2(_1844_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3502_ (.A1(_1698_),
    .A2(_1940_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3503_ (.A1(_1717_),
    .A2(net370),
    .B(_1936_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3504_ (.A1(_1812_),
    .A2(_0856_),
    .B1(_0857_),
    .B2(_1750_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _3505_ (.A1(_1698_),
    .A2(_1940_),
    .A3(_1938_),
    .B1(_0858_),
    .B2(net395),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3506_ (.A1(\minimax.regS_uc[14] ),
    .A2(_1786_),
    .B1(_0855_),
    .B2(_1831_),
    .C(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3507_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3508_ (.A1(_0854_),
    .A2(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3509_ (.A1(_0838_),
    .A2(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3510_ (.A1(_0853_),
    .A2(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3511_ (.A1(_0853_),
    .A2(_0863_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3512_ (.A1(_0758_),
    .A2(_0864_),
    .A3(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3513_ (.I(_0710_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3514_ (.I(_0854_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3515_ (.A1(_0868_),
    .A2(_0861_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3516_ (.I(_0703_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3517_ (.A1(_0271_),
    .A2(net7),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3518_ (.I(_0861_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3519_ (.A1(_0871_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3520_ (.A1(_0790_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3521_ (.A1(_0870_),
    .A2(_0873_),
    .B(_0874_),
    .C(_0844_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3522_ (.A1(net8),
    .A2(_0867_),
    .B1(_0869_),
    .B2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3523_ (.A1(_0583_),
    .A2(_0847_),
    .B(_0866_),
    .C(_0876_),
    .ZN(\minimax.aluX[14] ));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3524_ (.A1(_0606_),
    .A2(_0608_),
    .A3(_0610_),
    .B(_0238_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3525_ (.A1(\minimax.regS_ex[15] ),
    .A2(_0219_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3526_ (.A1(_0232_),
    .A2(_0825_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3527_ (.A1(_0187_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3528_ (.A1(\minimax.regS_uc[15] ),
    .A2(_0189_),
    .B1(_0878_),
    .B2(_0191_),
    .C(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3529_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3530_ (.A1(_0877_),
    .A2(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3531_ (.A1(_0648_),
    .A2(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3532_ (.I(_0883_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3533_ (.A1(_0648_),
    .A2(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3534_ (.A1(_0640_),
    .A2(_0871_),
    .A3(_0861_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3535_ (.A1(_0868_),
    .A2(_0872_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3536_ (.A1(_0849_),
    .A2(_0852_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3537_ (.A1(_0887_),
    .A2(_0888_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3538_ (.I(_0837_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3539_ (.A1(_0166_),
    .A2(_0891_),
    .A3(_0868_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3540_ (.I0(_0869_),
    .I1(_0892_),
    .S(_0889_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3541_ (.A1(_0166_),
    .A2(_0868_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3542_ (.A1(_0891_),
    .A2(_0868_),
    .A3(_0872_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3543_ (.A1(_0640_),
    .A2(_0891_),
    .A3(_0871_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3544_ (.A1(_0853_),
    .A2(_0894_),
    .B(_0895_),
    .C(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3545_ (.A1(_0890_),
    .A2(_0893_),
    .A3(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3546_ (.I0(_0884_),
    .I1(_0886_),
    .S(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3547_ (.A1(\bank1.rdata[15] ),
    .A2(_0511_),
    .B(_0740_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3548_ (.A1(_0877_),
    .A2(_0882_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3549_ (.A1(_0877_),
    .A2(_0882_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3550_ (.A1(_0680_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3551_ (.A1(_0870_),
    .A2(_0902_),
    .B(_0903_),
    .C(_0688_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3552_ (.A1(net9),
    .A2(_0718_),
    .B1(_0901_),
    .B2(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3553_ (.A1(_0591_),
    .A2(_0900_),
    .B(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3554_ (.A1(_0899_),
    .A2(_0906_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3555_ (.I(_0907_),
    .Z(\minimax.aluX[15] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3556_ (.A1(\bank1.rdata[16] ),
    .A2(_0739_),
    .B(_0716_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3557_ (.A1(_0891_),
    .A2(_0869_),
    .B1(_0862_),
    .B2(_0164_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3558_ (.A1(_0831_),
    .A2(_0837_),
    .A3(_0862_),
    .A4(_0883_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3559_ (.A1(_0638_),
    .A2(_0891_),
    .A3(_0873_),
    .A4(_0885_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3560_ (.A1(_0885_),
    .A2(_0909_),
    .B(_0910_),
    .C(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3561_ (.A1(_0287_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3562_ (.A1(_0837_),
    .A2(_0872_),
    .B(_0831_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3563_ (.A1(_0882_),
    .A2(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3564_ (.A1(_0871_),
    .A2(_0872_),
    .A3(_0901_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3565_ (.A1(_0721_),
    .A2(net8),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3566_ (.A1(_0917_),
    .A2(_0882_),
    .B(_0838_),
    .C(_0888_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3567_ (.A1(_0877_),
    .A2(_0915_),
    .B1(_0916_),
    .B2(_0838_),
    .C(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3568_ (.A1(_0822_),
    .A2(_0839_),
    .A3(_0912_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3569_ (.A1(_0919_),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3570_ (.A1(_0819_),
    .A2(_0848_),
    .A3(_0913_),
    .B(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3571_ (.A1(_0216_),
    .A2(_0835_),
    .A3(_0860_),
    .A4(_0881_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3572_ (.A1(_2049_),
    .A2(_0242_),
    .A3(_0244_),
    .A4(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3573_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3574_ (.I(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3575_ (.A1(_0651_),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3576_ (.A1(_0720_),
    .A2(net9),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3577_ (.I(_0219_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3578_ (.A1(\minimax.regS_ex[16] ),
    .A2(_0929_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3579_ (.A1(_1762_),
    .A2(_0825_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3580_ (.A1(_0188_),
    .A2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3581_ (.A1(\minimax.regS_uc[16] ),
    .A2(_0257_),
    .B1(_0930_),
    .B2(_0191_),
    .C(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3582_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3583_ (.A1(_0928_),
    .A2(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3584_ (.A1(_0927_),
    .A2(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3585_ (.A1(_0922_),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3586_ (.A1(_0695_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3587_ (.I(_0934_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3588_ (.A1(_0928_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3589_ (.A1(_0928_),
    .A2(_0939_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3590_ (.A1(_0782_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3591_ (.A1(_0697_),
    .A2(_0941_),
    .B(_0942_),
    .C(_0844_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3592_ (.A1(net10),
    .A2(_0867_),
    .B1(_0940_),
    .B2(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3593_ (.A1(_0374_),
    .A2(_0908_),
    .B(_0938_),
    .C(_0944_),
    .ZN(\minimax.aluX[16] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3594_ (.A1(\minimax.regS_ex[17] ),
    .A2(_0929_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3595_ (.A1(_1629_),
    .A2(_1631_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _3596_ (.A1(_1850_),
    .A2(_0856_),
    .A3(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3597_ (.A1(\minimax.regS_uc[17] ),
    .A2(_0189_),
    .B1(_0945_),
    .B2(_0191_),
    .C(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3598_ (.I(_0948_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3599_ (.I(_0288_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3600_ (.A1(_0950_),
    .A2(net10),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3601_ (.A1(_0949_),
    .A2(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3602_ (.A1(_0166_),
    .A2(_0928_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3603_ (.A1(_0922_),
    .A2(_0926_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3604_ (.A1(_0821_),
    .A2(net9),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3605_ (.A1(_0290_),
    .A2(_0934_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3606_ (.A1(_0955_),
    .A2(_0939_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3607_ (.A1(_0955_),
    .A2(_0956_),
    .B(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3608_ (.A1(_0815_),
    .A2(_0300_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3609_ (.A1(_0791_),
    .A2(_0324_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3610_ (.A1(_0791_),
    .A2(_0181_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3611_ (.I0(_0960_),
    .I1(_0961_),
    .S(_0177_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3612_ (.A1(_0213_),
    .A2(_0264_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3613_ (.A1(_0263_),
    .A2(_0265_),
    .B(_0959_),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3614_ (.A1(_0331_),
    .A2(_0332_),
    .A3(_0251_),
    .B(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3615_ (.A1(_0848_),
    .A2(_0913_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3616_ (.A1(_0919_),
    .A2(_0920_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3617_ (.A1(_0965_),
    .A2(_0966_),
    .B(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3618_ (.A1(_0968_),
    .A2(_0927_),
    .B(_0940_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3619_ (.A1(_0922_),
    .A2(_0953_),
    .B1(_0954_),
    .B2(_0958_),
    .C(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3620_ (.A1(_0952_),
    .A2(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3621_ (.A1(_0821_),
    .A2(net10),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3622_ (.A1(_0949_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3623_ (.A1(_0744_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3624_ (.A1(_0743_),
    .A2(_0973_),
    .B(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3625_ (.A1(_0949_),
    .A2(_0972_),
    .B1(_0975_),
    .B2(_0677_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3626_ (.A1(net11),
    .A2(_0799_),
    .B1(_0800_),
    .B2(_0971_),
    .C(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3627_ (.A1(_0400_),
    .A2(_0402_),
    .A3(_0798_),
    .B(_0977_),
    .ZN(\minimax.aluX[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3628_ (.I(_0710_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3629_ (.A1(_0926_),
    .A2(_0940_),
    .B1(_0935_),
    .B2(_0165_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3630_ (.I0(_0941_),
    .I1(_0935_),
    .S(_0926_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3631_ (.A1(_0639_),
    .A2(_0952_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3632_ (.A1(_0952_),
    .A2(_0979_),
    .B1(_0980_),
    .B2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3633_ (.I(_0924_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3634_ (.I(_0949_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3635_ (.A1(_0983_),
    .A2(_0955_),
    .B(_0984_),
    .C(_0956_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3636_ (.A1(_0983_),
    .A2(_0984_),
    .B(_0951_),
    .C(_0939_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3637_ (.A1(_0985_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3638_ (.A1(net10),
    .A2(_0934_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3639_ (.A1(_0928_),
    .A2(_0988_),
    .B(_0956_),
    .C(_0984_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3640_ (.A1(_0272_),
    .A2(_0835_),
    .A3(_0861_),
    .A4(_0881_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3641_ (.A1(_2027_),
    .A2(_0218_),
    .A3(_0229_),
    .A4(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3642_ (.A1(_0638_),
    .A2(_0991_),
    .A3(_0972_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3643_ (.A1(_0824_),
    .A2(_0983_),
    .A3(_0939_),
    .A4(_0949_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3644_ (.A1(_0955_),
    .A2(_0951_),
    .B1(_0989_),
    .B2(_0992_),
    .C(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3645_ (.A1(_0987_),
    .A2(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3646_ (.A1(_0968_),
    .A2(_0982_),
    .B(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3647_ (.A1(_0934_),
    .A2(_0948_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3648_ (.A1(_1850_),
    .A2(_0856_),
    .A3(_0946_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3649_ (.I(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3650_ (.I(\minimax.regS_ex[18] ),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3651_ (.I(\minimax.regS_uc[18] ),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3652_ (.I0(_1000_),
    .I1(_1001_),
    .S(_0189_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3653_ (.A1(_0999_),
    .A2(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3654_ (.A1(_0983_),
    .A2(_0997_),
    .B(_1003_),
    .C(_0164_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3655_ (.I(_0998_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3656_ (.A1(_1005_),
    .A2(_1002_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3657_ (.A1(_0990_),
    .A2(_0997_),
    .A3(_1003_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3658_ (.A1(_0638_),
    .A2(_1006_),
    .B1(_1007_),
    .B2(_0296_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3659_ (.A1(_0721_),
    .A2(net11),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3660_ (.A1(_1004_),
    .A2(_1008_),
    .B(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3661_ (.I(_0271_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3662_ (.A1(_1011_),
    .A2(net11),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3663_ (.A1(_1004_),
    .A2(_1008_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3664_ (.A1(_1012_),
    .A2(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3665_ (.A1(_1010_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3666_ (.A1(_0996_),
    .A2(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3667_ (.A1(_0812_),
    .A2(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_1009_),
    .A2(_1006_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3669_ (.I0(_0683_),
    .I1(_0744_),
    .S(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3670_ (.A1(_1012_),
    .A2(_1003_),
    .B1(_1019_),
    .B2(_0844_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3671_ (.A1(net12),
    .A2(_0978_),
    .B(_1017_),
    .C(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3672_ (.A1(_0417_),
    .A2(_0418_),
    .A3(_0798_),
    .B(_1021_),
    .ZN(\minimax.aluX[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3673_ (.I(_0812_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3674_ (.A1(_0933_),
    .A2(_0998_),
    .A3(_0948_),
    .A4(_1002_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3675_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3676_ (.A1(_0983_),
    .A2(_1024_),
    .B(_0824_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3677_ (.I(_0654_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3678_ (.A1(\minimax.regS_uc[19] ),
    .A2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3679_ (.I(_0179_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3680_ (.A1(\minimax.regS_ex[19] ),
    .A2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3681_ (.A1(_1005_),
    .A2(_1027_),
    .A3(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3682_ (.A1(_0950_),
    .A2(net12),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3683_ (.A1(_1030_),
    .A2(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3684_ (.I(_0947_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3685_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3686_ (.A1(\minimax.regS_uc[19] ),
    .A2(_0654_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3687_ (.A1(\minimax.regS_ex[19] ),
    .A2(_1028_),
    .B(_1034_),
    .C(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3688_ (.A1(_0821_),
    .A2(net12),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3689_ (.A1(_1036_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3690_ (.A1(_1032_),
    .A2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3691_ (.A1(_1025_),
    .A2(_1039_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3692_ (.A1(_1012_),
    .A2(_1013_),
    .B(_0968_),
    .C(_0982_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3693_ (.A1(_1012_),
    .A2(_1013_),
    .B(_0995_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3694_ (.A1(_1014_),
    .A2(_1041_),
    .A3(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3695_ (.A1(_1040_),
    .A2(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3696_ (.A1(_0790_),
    .A2(_1032_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3697_ (.A1(_0870_),
    .A2(_1032_),
    .B(_1045_),
    .C(_0688_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3698_ (.A1(net14),
    .A2(_0867_),
    .B1(_1038_),
    .B2(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3699_ (.I(_0740_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3700_ (.A1(net81),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3701_ (.A1(_1022_),
    .A2(_1044_),
    .B(_1047_),
    .C(_1049_),
    .ZN(\minimax.aluX[19] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3702_ (.A1(_0950_),
    .A2(net14),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3703_ (.A1(\minimax.regS_uc[20] ),
    .A2(_0190_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3704_ (.A1(\minimax.regS_ex[20] ),
    .A2(_0179_),
    .B(_1033_),
    .C(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3705_ (.I(_1052_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3706_ (.A1(_1050_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3707_ (.A1(_1050_),
    .A2(_1053_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3708_ (.I(_0998_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3709_ (.A1(_0933_),
    .A2(_1056_),
    .A3(_0948_),
    .A4(_1002_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3710_ (.A1(_1057_),
    .A2(_1036_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3711_ (.A1(_0925_),
    .A2(_1058_),
    .B(_0164_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3712_ (.A1(_1054_),
    .A2(_1055_),
    .B(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3713_ (.A1(_0950_),
    .A2(net14),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3714_ (.A1(_1061_),
    .A2(_1053_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3715_ (.A1(_1061_),
    .A2(_1052_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3716_ (.A1(_0926_),
    .A2(_1058_),
    .B1(_1062_),
    .B2(_1063_),
    .C(_0824_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3717_ (.A1(_1060_),
    .A2(_1064_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3718_ (.A1(_0982_),
    .A2(_1015_),
    .A3(_1040_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3719_ (.A1(_1024_),
    .A2(_1036_),
    .A3(_1031_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3720_ (.A1(_0164_),
    .A2(_1036_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3721_ (.A1(_0991_),
    .A2(_1067_),
    .B1(_1068_),
    .B2(_1037_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3722_ (.A1(_1025_),
    .A2(_1038_),
    .B(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3723_ (.A1(_0987_),
    .A2(_0994_),
    .A3(_1010_),
    .A4(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3724_ (.A1(_1009_),
    .A2(_1004_),
    .A3(_1008_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3725_ (.A1(_1024_),
    .A2(_1030_),
    .A3(_1037_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3726_ (.A1(_0824_),
    .A2(_1030_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3727_ (.A1(_0991_),
    .A2(_1073_),
    .B1(_1074_),
    .B2(_1031_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3728_ (.A1(_1025_),
    .A2(_1032_),
    .B1(_1070_),
    .B2(_1072_),
    .C(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3729_ (.A1(_1071_),
    .A2(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3730_ (.A1(_0968_),
    .A2(_1066_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3731_ (.A1(_1065_),
    .A2(_1078_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3732_ (.A1(_0694_),
    .A2(_1079_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3733_ (.I(_0686_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3734_ (.A1(_1081_),
    .A2(_1054_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3735_ (.A1(_0782_),
    .A2(_1054_),
    .B(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3736_ (.A1(_0781_),
    .A2(_1083_),
    .B(_1055_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3737_ (.A1(net15),
    .A2(_0978_),
    .B(_1080_),
    .C(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _3738_ (.A1(_0455_),
    .A2(_0456_),
    .A3(_0660_),
    .B(_1085_),
    .ZN(\minimax.aluX[20] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3739_ (.I(\minimax.regS_ex[21] ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3740_ (.I(\minimax.regS_uc[21] ),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _3741_ (.I0(_1086_),
    .I1(_1087_),
    .S(_0257_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3742_ (.A1(_1056_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3743_ (.A1(_0102_),
    .A2(_0990_),
    .A3(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3744_ (.A1(_1056_),
    .A2(_1088_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3745_ (.I(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3746_ (.A1(_0236_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3747_ (.A1(\minimax.regS_ex[19] ),
    .A2(\minimax.regS_ex[20] ),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3748_ (.A1(\minimax.regS_uc[19] ),
    .A2(\minimax.regS_uc[20] ),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3749_ (.I0(_1094_),
    .I1(_1095_),
    .S(_0826_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3750_ (.A1(_0096_),
    .A2(_0098_),
    .A3(_0228_),
    .A4(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3751_ (.A1(_0242_),
    .A2(_0999_),
    .A3(_1057_),
    .A4(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3752_ (.I0(_1090_),
    .I1(_1093_),
    .S(_1098_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3753_ (.I(_0110_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3754_ (.I(_1089_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3755_ (.A1(_0102_),
    .A2(_0990_),
    .B(_1101_),
    .C(_1100_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3756_ (.A1(_0720_),
    .A2(net15),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3757_ (.A1(_1100_),
    .A2(_1101_),
    .B(_1102_),
    .C(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3758_ (.A1(_0271_),
    .A2(net15),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3759_ (.A1(_0297_),
    .A2(_0923_),
    .A3(_1105_),
    .A4(_1092_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3760_ (.A1(_1100_),
    .A2(_1105_),
    .A3(_1101_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3761_ (.I0(_1106_),
    .I1(_1107_),
    .S(_1098_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3762_ (.A1(_1100_),
    .A2(_1101_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3763_ (.A1(_0236_),
    .A2(_1103_),
    .A3(_1092_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3764_ (.A1(_0297_),
    .A2(_0923_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3765_ (.A1(_1105_),
    .A2(_1109_),
    .B1(_1110_),
    .B2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3766_ (.A1(_1099_),
    .A2(_1104_),
    .B(_1108_),
    .C(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3767_ (.A1(_1059_),
    .A2(_1053_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3768_ (.A1(_1050_),
    .A2(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3769_ (.A1(_1065_),
    .A2(_1078_),
    .B(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3770_ (.A1(_1113_),
    .A2(_1116_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3771_ (.A1(_0695_),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(_1105_),
    .A2(_1101_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3773_ (.I0(_0792_),
    .I1(_1081_),
    .S(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3774_ (.A1(_1103_),
    .A2(_1092_),
    .B1(_1120_),
    .B2(_0801_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3775_ (.A1(net16),
    .A2(_0978_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3776_ (.A1(_0475_),
    .A2(_0767_),
    .B(_1118_),
    .C(_1122_),
    .ZN(\minimax.aluX[21] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3777_ (.A1(net85),
    .A2(_1048_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3778_ (.A1(_1099_),
    .A2(_1104_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3779_ (.I(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3780_ (.A1(_1108_),
    .A2(_1112_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3781_ (.A1(_1050_),
    .A2(_1052_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3782_ (.A1(_1061_),
    .A2(_1053_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3783_ (.I0(_1127_),
    .I1(_1128_),
    .S(_1059_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(_1126_),
    .A2(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3785_ (.A1(_1060_),
    .A2(_1064_),
    .B(_1113_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3786_ (.A1(_1125_),
    .A2(_1130_),
    .B1(_1131_),
    .B2(_1078_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3787_ (.I(\minimax.regS_ex[22] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3788_ (.A1(\minimax.regS_uc[22] ),
    .A2(_0654_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3789_ (.A1(_1133_),
    .A2(_0655_),
    .B(_0999_),
    .C(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3790_ (.A1(_0297_),
    .A2(_0923_),
    .A3(_1092_),
    .A4(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3791_ (.A1(\minimax.regS_uc[22] ),
    .A2(_0826_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3792_ (.A1(\minimax.regS_ex[22] ),
    .A2(_1028_),
    .B(_1033_),
    .C(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3793_ (.A1(_1100_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3794_ (.I0(_1136_),
    .I1(_1139_),
    .S(_1098_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3795_ (.A1(_0236_),
    .A2(_1135_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3796_ (.A1(_0110_),
    .A2(_1138_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3797_ (.A1(_1093_),
    .A2(_1138_),
    .B1(_1141_),
    .B2(_1111_),
    .C(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3798_ (.A1(_0821_),
    .A2(net16),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3799_ (.A1(_1140_),
    .A2(_1143_),
    .B(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3800_ (.A1(_1144_),
    .A2(_1140_),
    .A3(_1143_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3801_ (.A1(_1145_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3802_ (.A1(_1132_),
    .A2(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3803_ (.A1(_1011_),
    .A2(net16),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3804_ (.A1(_1144_),
    .A2(_1135_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3805_ (.I0(_0792_),
    .I1(_0697_),
    .S(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3806_ (.A1(_1149_),
    .A2(_1138_),
    .B1(_1151_),
    .B2(_0781_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3807_ (.A1(net17),
    .A2(_0780_),
    .B1(_0758_),
    .B2(_1148_),
    .C(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3808_ (.A1(_1123_),
    .A2(_1153_),
    .ZN(\minimax.aluX[22] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3809_ (.A1(\minimax.regS_ex[22] ),
    .A2(_1094_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3810_ (.A1(\minimax.regS_uc[22] ),
    .A2(_1095_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3811_ (.I0(_1154_),
    .I1(_1155_),
    .S(_0190_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(_1091_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3813_ (.A1(_0924_),
    .A2(_1024_),
    .A3(_1157_),
    .B(_0163_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3814_ (.A1(\minimax.regS_ex[23] ),
    .A2(_0947_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3815_ (.A1(\minimax.regS_uc[23] ),
    .A2(_0947_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3816_ (.I0(_1159_),
    .I1(_1160_),
    .S(_0190_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3817_ (.I(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3818_ (.A1(_0720_),
    .A2(net17),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_4 _3819_ (.A1(_1158_),
    .A2(_1162_),
    .A3(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3820_ (.A1(_0812_),
    .A2(_1146_),
    .A3(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3821_ (.A1(_1132_),
    .A2(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3822_ (.A1(_1140_),
    .A2(_1143_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3823_ (.A1(_1149_),
    .A2(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3824_ (.A1(_1125_),
    .A2(_1130_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3825_ (.A1(_1169_),
    .A2(_1167_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3826_ (.A1(_1169_),
    .A2(_1167_),
    .B(_1149_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3827_ (.A1(_1164_),
    .A2(_1170_),
    .A3(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3828_ (.A1(_1078_),
    .A2(_1131_),
    .A3(_1168_),
    .A4(_1164_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3829_ (.A1(_1168_),
    .A2(_1164_),
    .B(_1172_),
    .C(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3830_ (.I(_1163_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3831_ (.A1(_1162_),
    .A2(_1175_),
    .B(_0696_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3832_ (.A1(_0743_),
    .A2(_1162_),
    .A3(_1175_),
    .B(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3833_ (.A1(_1162_),
    .A2(_1175_),
    .B1(_1177_),
    .B2(_0719_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3834_ (.A1(net18),
    .A2(_0799_),
    .B1(_0800_),
    .B2(_1174_),
    .C(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3835_ (.A1(_0501_),
    .A2(_0767_),
    .B(_1166_),
    .C(_1179_),
    .ZN(\minimax.aluX[23] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3836_ (.A1(net87),
    .A2(_1048_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3837_ (.A1(_0982_),
    .A2(_1010_),
    .A3(_1014_),
    .A4(_1040_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3838_ (.A1(_1145_),
    .A2(_1146_),
    .A3(_1164_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3839_ (.A1(_1131_),
    .A2(_1182_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3840_ (.A1(_1181_),
    .A2(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3841_ (.A1(_1158_),
    .A2(_1162_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3842_ (.A1(_1175_),
    .A2(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3843_ (.A1(_1126_),
    .A2(_1129_),
    .B1(_1149_),
    .B2(_1167_),
    .C(_1124_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3844_ (.A1(_1175_),
    .A2(_1185_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3845_ (.A1(_1146_),
    .A2(_1186_),
    .A3(_1187_),
    .B(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3846_ (.A1(_1071_),
    .A2(_1076_),
    .B(_1131_),
    .C(_1182_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3847_ (.A1(_1189_),
    .A2(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3848_ (.A1(_0968_),
    .A2(_1184_),
    .B(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3849_ (.A1(\minimax.regS_uc[24] ),
    .A2(_0826_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3850_ (.A1(\minimax.regS_ex[24] ),
    .A2(_0657_),
    .A3(_0929_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3851_ (.A1(_1056_),
    .A2(_1193_),
    .A3(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3852_ (.I(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3853_ (.A1(_0721_),
    .A2(net18),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3854_ (.A1(_1196_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3855_ (.A1(_0999_),
    .A2(_1193_),
    .A3(_1194_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3856_ (.I(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3857_ (.A1(_0950_),
    .A2(net18),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3858_ (.A1(_1200_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3859_ (.A1(_1198_),
    .A2(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3860_ (.A1(_1056_),
    .A2(_1088_),
    .A3(_1156_),
    .A4(_1161_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3861_ (.A1(_1023_),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3862_ (.A1(_0991_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3863_ (.I(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3864_ (.A1(_0166_),
    .A2(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3865_ (.A1(_1203_),
    .A2(_1208_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3866_ (.A1(_1192_),
    .A2(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3867_ (.A1(_0695_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3868_ (.A1(_0790_),
    .A2(_1202_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3869_ (.A1(_0870_),
    .A2(_1202_),
    .B(_1212_),
    .C(_0688_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3870_ (.A1(net19),
    .A2(_0780_),
    .B1(_1198_),
    .B2(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3871_ (.A1(_1180_),
    .A2(_1211_),
    .A3(_1214_),
    .ZN(\minimax.aluX[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3872_ (.A1(_0721_),
    .A2(net19),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3873_ (.I(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3874_ (.A1(\minimax.regS_uc[25] ),
    .A2(_1026_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3875_ (.A1(\minimax.regS_ex[25] ),
    .A2(_0699_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3876_ (.A1(_1005_),
    .A2(_1217_),
    .A3(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3877_ (.A1(_1216_),
    .A2(_1219_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3878_ (.A1(_1216_),
    .A2(_1219_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3879_ (.A1(_1220_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3880_ (.A1(_1181_),
    .A2(_1183_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3881_ (.A1(_1189_),
    .A2(_1190_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3882_ (.A1(_0922_),
    .A2(_1223_),
    .B(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3883_ (.A1(_1196_),
    .A2(_1201_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3884_ (.A1(_1195_),
    .A2(_1201_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3885_ (.A1(_1225_),
    .A2(_1226_),
    .B(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3886_ (.A1(_1207_),
    .A2(_1192_),
    .A3(_1198_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3887_ (.A1(_1200_),
    .A2(_1201_),
    .B(_0640_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3888_ (.A1(_0640_),
    .A2(_1228_),
    .B1(_1229_),
    .B2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3889_ (.A1(_1222_),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3890_ (.A1(_0681_),
    .A2(_1221_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3891_ (.A1(_0870_),
    .A2(_1221_),
    .B(_1233_),
    .C(_0677_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3892_ (.A1(net20),
    .A2(_0867_),
    .B1(_1220_),
    .B2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3893_ (.A1(net88),
    .A2(_0741_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3894_ (.A1(_1022_),
    .A2(_1232_),
    .B(_1235_),
    .C(_1236_),
    .ZN(\minimax.aluX[25] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3895_ (.A1(_1206_),
    .A2(_1201_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3896_ (.A1(_0991_),
    .A2(_1205_),
    .B(_1200_),
    .C(_1197_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3897_ (.A1(_1200_),
    .A2(_1237_),
    .B(_1238_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3898_ (.A1(_1207_),
    .A2(_1198_),
    .B1(_1203_),
    .B2(_0651_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3899_ (.A1(_1222_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3900_ (.A1(_0236_),
    .A2(_1222_),
    .A3(_1239_),
    .B(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3901_ (.A1(_1206_),
    .A2(_1199_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3902_ (.A1(_1200_),
    .A2(_1215_),
    .B1(_1243_),
    .B2(_0165_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3903_ (.A1(_0639_),
    .A2(_1196_),
    .A3(_1219_),
    .B(_1216_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3904_ (.A1(_1196_),
    .A2(_1215_),
    .B1(_1227_),
    .B2(_0639_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3905_ (.A1(_1207_),
    .A2(_1198_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3906_ (.A1(_1207_),
    .A2(_1196_),
    .A3(_1216_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3907_ (.A1(_1197_),
    .A2(_1245_),
    .B1(_1247_),
    .B2(_1219_),
    .C(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3908_ (.A1(_1219_),
    .A2(_1244_),
    .B(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3909_ (.I(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3910_ (.A1(_1192_),
    .A2(_1242_),
    .B(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3911_ (.A1(_1011_),
    .A2(net20),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3912_ (.A1(\minimax.regS_uc[26] ),
    .A2(_0655_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3913_ (.A1(\minimax.regS_ex[26] ),
    .A2(_1028_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3914_ (.A1(_1005_),
    .A2(_1254_),
    .A3(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3915_ (.I(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _3916_ (.A1(_1024_),
    .A2(_1204_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3917_ (.A1(\minimax.regS_ex[24] ),
    .A2(\minimax.regS_ex[25] ),
    .A3(_0654_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3918_ (.A1(\minimax.regS_uc[24] ),
    .A2(\minimax.regS_uc[25] ),
    .A3(_1028_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3919_ (.A1(_1259_),
    .A2(_1260_),
    .B(_1005_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3920_ (.A1(_0925_),
    .A2(_1258_),
    .A3(_1261_),
    .B(_0831_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3921_ (.A1(_1257_),
    .A2(_1262_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3922_ (.A1(_1253_),
    .A2(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3923_ (.A1(_1252_),
    .A2(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3924_ (.A1(_0722_),
    .A2(net20),
    .A3(_1256_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3925_ (.I0(_0683_),
    .I1(_1081_),
    .S(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3926_ (.A1(_1257_),
    .A2(_1253_),
    .B1(_1267_),
    .B2(_0801_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3927_ (.A1(net21),
    .A2(_0978_),
    .B(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3928_ (.A1(_0542_),
    .A2(_0767_),
    .B1(_1265_),
    .B2(_0649_),
    .C(_1269_),
    .ZN(\minimax.aluX[26] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3929_ (.A1(_1253_),
    .A2(_1263_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3930_ (.A1(_1011_),
    .A2(net21),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3931_ (.A1(\minimax.regS_uc[27] ),
    .A2(_0257_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3932_ (.A1(\minimax.regS_ex[27] ),
    .A2(_0179_),
    .B(_0947_),
    .C(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3933_ (.I(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3934_ (.A1(\minimax.regS_ex[25] ),
    .A2(\minimax.regS_ex[26] ),
    .A3(_1033_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3935_ (.A1(\minimax.regS_uc[25] ),
    .A2(\minimax.regS_uc[26] ),
    .A3(_1033_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3936_ (.I0(_1275_),
    .I1(_1276_),
    .S(_0826_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3937_ (.A1(_0999_),
    .A2(_1193_),
    .A3(_1194_),
    .A4(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3938_ (.A1(_0925_),
    .A2(_1258_),
    .A3(_1274_),
    .A4(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3939_ (.A1(_0163_),
    .A2(_0924_),
    .A3(_1273_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3940_ (.A1(_0163_),
    .A2(_1258_),
    .A3(_1273_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3941_ (.A1(_0163_),
    .A2(_1273_),
    .A3(_1278_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3942_ (.A1(_0831_),
    .A2(_1274_),
    .B(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _3943_ (.A1(_1279_),
    .A2(_1280_),
    .A3(_1281_),
    .A4(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3944_ (.A1(_1271_),
    .A2(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3945_ (.A1(_1270_),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3946_ (.A1(_1253_),
    .A2(_1263_),
    .B(_1252_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3947_ (.I0(_1286_),
    .I1(_1285_),
    .S(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3948_ (.A1(net90),
    .A2(_1048_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3949_ (.A1(_1270_),
    .A2(_1285_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3950_ (.I(_1271_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3951_ (.A1(_1291_),
    .A2(_1274_),
    .B(_0696_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3952_ (.A1(_0743_),
    .A2(_1291_),
    .A3(_1274_),
    .B(_1292_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3953_ (.A1(_1291_),
    .A2(_1274_),
    .B1(_1293_),
    .B2(_0777_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _3954_ (.A1(net22),
    .A2(_0799_),
    .B1(_0800_),
    .B2(_1290_),
    .C(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3955_ (.A1(_1022_),
    .A2(_1288_),
    .B(_1289_),
    .C(_1295_),
    .ZN(\minimax.aluX[27] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3956_ (.I(_1242_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3957_ (.A1(_1264_),
    .A2(_1285_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3958_ (.A1(_1250_),
    .A2(_1263_),
    .B(_1253_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3959_ (.A1(_1250_),
    .A2(_1263_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3960_ (.A1(_1291_),
    .A2(_1284_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3961_ (.A1(_1298_),
    .A2(_1299_),
    .B(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3962_ (.A1(_1291_),
    .A2(_1284_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3963_ (.A1(_1225_),
    .A2(_1296_),
    .A3(_1297_),
    .B1(_1301_),
    .B2(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3964_ (.A1(_0722_),
    .A2(net22),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _3965_ (.I0(\minimax.regS_ex[28] ),
    .I1(\minimax.regS_uc[28] ),
    .S(_0655_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3966_ (.A1(_1034_),
    .A2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3967_ (.A1(_1195_),
    .A2(_1273_),
    .A3(_1277_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3968_ (.A1(_1206_),
    .A2(_1307_),
    .B(_0165_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3969_ (.A1(_1306_),
    .A2(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3970_ (.A1(_1304_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3971_ (.A1(_1304_),
    .A2(_1309_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3972_ (.A1(_1310_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3973_ (.A1(_1303_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3974_ (.A1(_1304_),
    .A2(_1306_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3975_ (.A1(_1081_),
    .A2(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3976_ (.A1(_0782_),
    .A2(_1314_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3977_ (.A1(_1304_),
    .A2(_1306_),
    .B1(_1316_),
    .B2(_0844_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3978_ (.A1(net23),
    .A2(_0867_),
    .B(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _3979_ (.A1(_0565_),
    .A2(_0767_),
    .B1(_1313_),
    .B2(_0812_),
    .C(_1318_),
    .ZN(\minimax.aluX[28] ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3980_ (.A1(_1296_),
    .A2(_1297_),
    .A3(_1310_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3981_ (.A1(_1271_),
    .A2(_1284_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3982_ (.A1(_1271_),
    .A2(_1284_),
    .B(_1270_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3983_ (.A1(_1320_),
    .A2(_1321_),
    .B(_1311_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3984_ (.A1(_1250_),
    .A2(_1297_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3985_ (.A1(_1322_),
    .A2(_1323_),
    .B(_1310_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3986_ (.A1(_1192_),
    .A2(_1319_),
    .B(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3987_ (.A1(_0722_),
    .A2(net23),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3988_ (.A1(\minimax.regS_uc[29] ),
    .A2(_0655_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3989_ (.A1(\minimax.regS_ex[29] ),
    .A2(_0699_),
    .B(_1034_),
    .C(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3990_ (.A1(_0925_),
    .A2(_1258_),
    .A3(_1305_),
    .A4(_1307_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3991_ (.A1(_0638_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3992_ (.A1(_1328_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3993_ (.A1(_1326_),
    .A2(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3994_ (.A1(_1326_),
    .A2(_1331_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3995_ (.I(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3996_ (.A1(_1332_),
    .A2(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3997_ (.A1(_1325_),
    .A2(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3998_ (.A1(net92),
    .A2(_1048_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3999_ (.A1(_1326_),
    .A2(_1328_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4000_ (.A1(_1081_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4001_ (.A1(_0782_),
    .A2(_1338_),
    .B(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4002_ (.A1(_1326_),
    .A2(_1328_),
    .B1(_1340_),
    .B2(_0801_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4003_ (.A1(net25),
    .A2(_0978_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4004_ (.A1(_1022_),
    .A2(_1336_),
    .B(_1337_),
    .C(_1342_),
    .ZN(\minimax.aluX[29] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4005_ (.A1(_0722_),
    .A2(net25),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4006_ (.I0(\minimax.regS_ex[30] ),
    .I1(\minimax.regS_uc[30] ),
    .S(_1026_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4007_ (.A1(_1034_),
    .A2(_1344_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4008_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4009_ (.A1(_0651_),
    .A2(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4010_ (.A1(_1345_),
    .A2(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4011_ (.A1(_1343_),
    .A2(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4012_ (.A1(_1343_),
    .A2(_1348_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4013_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4014_ (.A1(_1334_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4015_ (.A1(_1325_),
    .A2(_1332_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4016_ (.A1(_1325_),
    .A2(_1352_),
    .B1(_1353_),
    .B2(_1351_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4017_ (.I(_1332_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_1334_),
    .A2(_1351_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4019_ (.A1(_1355_),
    .A2(_1351_),
    .B(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4020_ (.A1(_1343_),
    .A2(_1345_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4021_ (.I0(_0683_),
    .I1(_0744_),
    .S(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4022_ (.A1(_1343_),
    .A2(_1345_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4023_ (.A1(_0688_),
    .A2(_1359_),
    .B(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4024_ (.A1(net26),
    .A2(_0664_),
    .B1(_0694_),
    .B2(_1357_),
    .C(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4025_ (.A1(net94),
    .A2(_0741_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4026_ (.A1(_1022_),
    .A2(_1354_),
    .B(_1362_),
    .C(_1363_),
    .ZN(\minimax.aluX[30] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4027_ (.A1(_1011_),
    .A2(net26),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4028_ (.A1(\minimax.regS_uc[31] ),
    .A2(_1026_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4029_ (.A1(\minimax.regS_ex[31] ),
    .A2(_0699_),
    .B(_1034_),
    .C(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4030_ (.A1(_1344_),
    .A2(_1346_),
    .B(_0651_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4031_ (.A1(_1364_),
    .A2(_1366_),
    .A3(_1367_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4032_ (.I(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4033_ (.A1(_1343_),
    .A2(_1348_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4034_ (.A1(_1325_),
    .A2(_1370_),
    .B(_1350_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4035_ (.A1(_1350_),
    .A2(_1368_),
    .B(_1333_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4036_ (.A1(_1192_),
    .A2(_1319_),
    .B(_1372_),
    .C(_1324_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4037_ (.A1(_1325_),
    .A2(_1355_),
    .B1(_1349_),
    .B2(_1369_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4038_ (.A1(_1369_),
    .A2(_1371_),
    .B(_1373_),
    .C(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4039_ (.I(_1350_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4040_ (.A1(_1334_),
    .A2(_1349_),
    .B1(_1376_),
    .B2(_1332_),
    .C(_1369_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4041_ (.A1(_1334_),
    .A2(_1370_),
    .B1(_1350_),
    .B2(_1332_),
    .C(_1368_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4042_ (.A1(_1377_),
    .A2(_1378_),
    .B(_0694_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4043_ (.A1(_0130_),
    .A2(_0710_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4044_ (.A1(_1366_),
    .A2(_1380_),
    .B(_1364_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4045_ (.A1(_1364_),
    .A2(_1366_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4046_ (.A1(_0792_),
    .A2(_1382_),
    .A3(_1380_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4047_ (.A1(_0790_),
    .A2(_1381_),
    .B(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4048_ (.A1(_1364_),
    .A2(_1366_),
    .B1(_1384_),
    .B2(_0781_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4049_ (.I(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4050_ (.A1(_0599_),
    .A2(_0661_),
    .B1(_1375_),
    .B2(_1379_),
    .C(_1386_),
    .ZN(\minimax.aluX[31] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _4051_ (.I(_0670_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4052_ (.A1(_0662_),
    .A2(_0641_),
    .B(_0725_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4053_ (.A1(_0648_),
    .A2(_0730_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4054_ (.A1(_1771_),
    .A2(_1388_),
    .B(_1389_),
    .C(_0740_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4055_ (.A1(_1387_),
    .A2(_1390_),
    .B(_1743_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4056_ (.A1(_1387_),
    .A2(_1390_),
    .B(_2034_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4057_ (.I(\minimax.dly16_slli_setrs ),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4058_ (.I(\minimax.dly16_slli_setrs ),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(_1392_),
    .A2(_0673_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4060_ (.A1(_0671_),
    .A2(_0642_),
    .B(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4061_ (.A1(_0109_),
    .A2(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4062_ (.I(\minimax.inst[7] ),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4063_ (.A1(_1629_),
    .A2(_1679_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4064_ (.A1(_1665_),
    .A2(_1397_),
    .B(_1847_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4065_ (.I(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4066_ (.A1(_1649_),
    .A2(_0668_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4067_ (.A1(net408),
    .A2(_1722_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4068_ (.A1(_1400_),
    .A2(_0672_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _4069_ (.I(_1402_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4070_ (.A1(_0641_),
    .A2(net408),
    .B(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _4071_ (.A1(_1399_),
    .A2(_1404_),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _4072_ (.A1(_1391_),
    .A2(\minimax.dra[0] ),
    .B1(_1395_),
    .B2(_1646_),
    .C1(_1396_),
    .C2(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4073_ (.I(_1406_),
    .ZN(\minimax.addrS_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4074_ (.A1(\minimax.op16_lwsp ),
    .A2(_1925_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4075_ (.A1(_1391_),
    .A2(\minimax.dra[1] ),
    .B1(_1395_),
    .B2(_1643_),
    .C(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(_2043_),
    .A2(_1405_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4077_ (.A1(_1408_),
    .A2(_1409_),
    .ZN(\minimax.addrS_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _4078_ (.A1(_1391_),
    .A2(\minimax.dra[2] ),
    .B1(_1395_),
    .B2(_0698_),
    .C1(_1815_),
    .C2(_1405_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4079_ (.I(_1410_),
    .ZN(\minimax.addrS_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4080_ (.A1(_0662_),
    .A2(_1771_),
    .B(_1404_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4081_ (.A1(_1391_),
    .A2(\minimax.dra[3] ),
    .B1(_1394_),
    .B2(_0674_),
    .C(_1399_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4082_ (.A1(_0195_),
    .A2(_1411_),
    .B(_1412_),
    .ZN(\minimax.addrS_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4083_ (.A1(_0233_),
    .A2(_1394_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4084_ (.A1(_1391_),
    .A2(\minimax.dra[4] ),
    .B1(_1404_),
    .B2(_0662_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _4085_ (.A1(_1413_),
    .A2(_1414_),
    .ZN(\minimax.addrS_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4086_ (.A1(\minimax.dly16_slli_setrd ),
    .A2(_1650_),
    .A3(_0671_),
    .A4(_0672_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4087_ (.A1(net364),
    .A2(_0646_),
    .A3(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _4088_ (.A1(\minimax.dly16_slli_setrd ),
    .A2(_0740_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4089_ (.A1(_0233_),
    .A2(_1814_),
    .B1(_1417_),
    .B2(\minimax.dra[4] ),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4090_ (.A1(_1848_),
    .A2(_1416_),
    .B(_1418_),
    .ZN(\minimax.addrD_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4091_ (.A1(_1702_),
    .A2(_1696_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4092_ (.A1(_1640_),
    .A2(_1419_),
    .B(_1626_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4093_ (.A1(_1646_),
    .A2(\minimax.op16_lw ),
    .B1(_1420_),
    .B2(_1396_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4094_ (.I(_1701_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4095_ (.A1(_1422_),
    .A2(net2),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4096_ (.A1(_1421_),
    .A2(_1423_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4097_ (.A1(_1643_),
    .A2(\minimax.op16_lw ),
    .B1(_1420_),
    .B2(_2043_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_1422_),
    .A2(net13),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_1424_),
    .A2(_1425_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4100_ (.A1(_0698_),
    .A2(\minimax.op16_lw ),
    .B1(_1420_),
    .B2(_1815_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_1422_),
    .A2(net24),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4102_ (.A1(_1426_),
    .A2(_1427_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4103_ (.A1(_1422_),
    .A2(net27),
    .B1(_1420_),
    .B2(_0130_),
    .C(\minimax.op16_lw ),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4104_ (.I(_1428_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4105_ (.A1(_1422_),
    .A2(net28),
    .B1(_1420_),
    .B2(_0662_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4106_ (.I(_1429_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4107_ (.A1(_1725_),
    .A2(_0657_),
    .B(_1401_),
    .C(_1961_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4108_ (.I(_1748_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4109_ (.A1(_2033_),
    .A2(net393),
    .A3(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4110_ (.I(_1431_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4111_ (.I(_1723_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4112_ (.I(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4113_ (.A1(\minimax.regS_ex[11] ),
    .A2(\minimax.regS_ex[14] ),
    .A3(\minimax.regS_ex[15] ),
    .A4(\minimax.regS_ex[16] ),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4114_ (.A1(\minimax.regS_ex[17] ),
    .A2(\minimax.regS_ex[18] ),
    .A3(\minimax.regS_ex[21] ),
    .A4(\minimax.regS_ex[23] ),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4115_ (.A1(\minimax.regS_ex[12] ),
    .A2(\minimax.regS_ex[13] ),
    .A3(\minimax.regS_ex[25] ),
    .A4(\minimax.regS_ex[26] ),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4116_ (.A1(_0220_),
    .A2(_1434_),
    .A3(_1435_),
    .A4(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4117_ (.A1(\minimax.regS_ex[5] ),
    .A2(\minimax.regS_ex[6] ),
    .A3(\minimax.regS_ex[7] ),
    .A4(\minimax.regS_ex[8] ),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4118_ (.A1(\minimax.regS_ex[24] ),
    .A2(\minimax.regS_ex[27] ),
    .A3(\minimax.regS_ex[28] ),
    .A4(\minimax.regS_ex[29] ),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4119_ (.A1(\minimax.regS_ex[4] ),
    .A2(\minimax.regS_ex[30] ),
    .A3(\minimax.regS_ex[31] ),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4120_ (.A1(_1154_),
    .A2(_1438_),
    .A3(_1439_),
    .A4(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4121_ (.A1(_1952_),
    .A2(_1437_),
    .A3(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4122_ (.A1(\minimax.regS_uc[12] ),
    .A2(\minimax.regS_uc[13] ),
    .A3(\minimax.regS_uc[25] ),
    .A4(\minimax.regS_uc[26] ),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4123_ (.A1(\minimax.regS_uc[15] ),
    .A2(\minimax.regS_uc[17] ),
    .A3(\minimax.regS_uc[18] ),
    .A4(\minimax.regS_uc[21] ),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4124_ (.A1(\minimax.regS_uc[11] ),
    .A2(\minimax.regS_uc[14] ),
    .A3(\minimax.regS_uc[16] ),
    .A4(\minimax.regS_uc[23] ),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4125_ (.A1(_0223_),
    .A2(_1443_),
    .A3(_1444_),
    .A4(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4126_ (.A1(\minimax.regS_uc[5] ),
    .A2(\minimax.regS_uc[6] ),
    .A3(\minimax.regS_uc[7] ),
    .A4(\minimax.regS_uc[8] ),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4127_ (.A1(\minimax.regS_uc[24] ),
    .A2(\minimax.regS_uc[27] ),
    .A3(\minimax.regS_uc[28] ),
    .A4(\minimax.regS_uc[29] ),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4128_ (.A1(\minimax.regS_uc[4] ),
    .A2(\minimax.regS_uc[30] ),
    .A3(\minimax.regS_uc[31] ),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4129_ (.A1(_1155_),
    .A2(_1447_),
    .A3(_1448_),
    .A4(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4130_ (.A1(_1946_),
    .A2(_1446_),
    .A3(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4131_ (.I0(_1442_),
    .I1(_1451_),
    .S(_0084_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4132_ (.A1(_1812_),
    .A2(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4133_ (.A1(_1847_),
    .A2(_1665_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4134_ (.A1(_1453_),
    .A2(_1454_),
    .B(_0665_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4135_ (.I(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4136_ (.I(_1456_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4137_ (.I(_1457_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4138_ (.A1(_1961_),
    .A2(_1433_),
    .A3(_1742_),
    .A4(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4139_ (.I(_1459_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4140_ (.A1(\minimax.regS_uc[1] ),
    .A2(_0656_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4141_ (.A1(_1863_),
    .A2(_0656_),
    .B(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(_1433_),
    .A2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(\minimax.pc_execute[1] ),
    .A2(_1403_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4144_ (.A1(_1658_),
    .A2(_1463_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4145_ (.A1(\minimax.pc_fetch[1] ),
    .A2(_1634_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4146_ (.A1(_1433_),
    .A2(_1742_),
    .A3(_1458_),
    .A4(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4147_ (.A1(_1458_),
    .A2(_1464_),
    .B(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4148_ (.A1(_1462_),
    .A2(_1467_),
    .B(_2033_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4149_ (.I(_1961_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4150_ (.A1(_1432_),
    .A2(_1742_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4151_ (.A1(\minimax.pc_fetch[1] ),
    .A2(_1639_),
    .A3(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4152_ (.A1(_1643_),
    .A2(\minimax.pc_execute[1] ),
    .A3(_1456_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4153_ (.A1(_1458_),
    .A2(_1470_),
    .B(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4154_ (.A1(_1811_),
    .A2(\minimax.pc_execute[2] ),
    .A3(_1402_),
    .A4(_1456_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(\minimax.pc_fetch[2] ),
    .A2(_0657_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4156_ (.I(\minimax.pc_execute[2] ),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4157_ (.I0(_1474_),
    .I1(_1475_),
    .S(_1455_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4158_ (.A1(_1432_),
    .A2(_0701_),
    .B1(_1456_),
    .B2(_0698_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4159_ (.A1(_1432_),
    .A2(_1476_),
    .B(_1477_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_1473_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4161_ (.A1(_1472_),
    .A2(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4162_ (.A1(_1468_),
    .A2(_1480_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4163_ (.I(_1455_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4164_ (.A1(_1481_),
    .A2(_1470_),
    .B(_1471_),
    .C(_1473_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4165_ (.A1(_1478_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4166_ (.A1(_1940_),
    .A2(_0946_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4167_ (.A1(_1453_),
    .A2(_1454_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4168_ (.A1(\minimax.regS_ex[3] ),
    .A2(_0929_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4169_ (.A1(\minimax.regS_uc[3] ),
    .A2(_0178_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4170_ (.A1(_1486_),
    .A2(_1487_),
    .B(_1402_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4171_ (.A1(_0232_),
    .A2(_1484_),
    .B1(_1485_),
    .B2(_0130_),
    .C(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4172_ (.A1(\minimax.pc_fetch[3] ),
    .A2(_1469_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4173_ (.I(\minimax.pc_execute[3] ),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4174_ (.I0(_1490_),
    .I1(_1491_),
    .S(_1455_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4175_ (.A1(_1483_),
    .A2(_1489_),
    .A3(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4176_ (.A1(_1468_),
    .A2(_1493_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(\minimax.pc_fetch[4] ),
    .A2(_1469_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4178_ (.A1(_1456_),
    .A2(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4179_ (.A1(\minimax.pc_execute[4] ),
    .A2(_1481_),
    .B(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4180_ (.I0(\minimax.regS_ex[4] ),
    .I1(\minimax.regS_uc[4] ),
    .S(_1026_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4181_ (.A1(_1432_),
    .A2(_1497_),
    .B1(_1481_),
    .B2(_0234_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4182_ (.A1(_1496_),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(_1489_),
    .A2(_1492_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4184_ (.A1(_1478_),
    .A2(_1482_),
    .A3(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4185_ (.A1(_1489_),
    .A2(_1492_),
    .B(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4186_ (.A1(_1499_),
    .A2(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4187_ (.A1(_1468_),
    .A2(_1503_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4188_ (.I(_1455_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4189_ (.I(_1469_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4190_ (.A1(\minimax.pc_fetch[5] ),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(\minimax.pc_execute[5] ),
    .A2(_1504_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4192_ (.A1(_1504_),
    .A2(_1506_),
    .B(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4193_ (.A1(_1645_),
    .A2(_1481_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4194_ (.A1(_1403_),
    .A2(_1973_),
    .B(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4195_ (.A1(_1508_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4196_ (.I(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_1508_),
    .A2(_1510_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_1512_),
    .A2(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4199_ (.A1(_1496_),
    .A2(_1498_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4200_ (.A1(_1496_),
    .A2(_1498_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4201_ (.A1(_1515_),
    .A2(_1502_),
    .B(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4202_ (.A1(_1514_),
    .A2(_1517_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4203_ (.A1(_1468_),
    .A2(_1518_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4204_ (.A1(_1511_),
    .A2(_1517_),
    .B(_1513_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4205_ (.A1(\minimax.regS_ex[6] ),
    .A2(_0929_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4206_ (.A1(\minimax.regS_uc[6] ),
    .A2(_0178_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4207_ (.A1(_1520_),
    .A2(_1521_),
    .B(_1403_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4208_ (.A1(_1396_),
    .A2(_1484_),
    .B1(_1485_),
    .B2(_0674_),
    .C(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(\minimax.pc_fetch[6] ),
    .A2(_1505_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4210_ (.A1(_1504_),
    .A2(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4211_ (.A1(\minimax.pc_execute[6] ),
    .A2(_1457_),
    .B(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4212_ (.A1(_1523_),
    .A2(_1526_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4213_ (.A1(_1523_),
    .A2(_1526_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4214_ (.A1(_1527_),
    .A2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4215_ (.A1(_1519_),
    .A2(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4216_ (.A1(_1468_),
    .A2(_1530_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4217_ (.I(_1876_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4218_ (.I(_1527_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4219_ (.A1(_1519_),
    .A2(_1532_),
    .B(_1528_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4220_ (.A1(\minimax.regS_uc[7] ),
    .A2(_0656_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4221_ (.A1(_2052_),
    .A2(_0656_),
    .B(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4222_ (.A1(_0233_),
    .A2(_1504_),
    .B1(_1535_),
    .B2(_1433_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4223_ (.A1(\minimax.pc_fetch[7] ),
    .A2(_1505_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4224_ (.A1(_1481_),
    .A2(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4225_ (.A1(\minimax.pc_execute[7] ),
    .A2(_1457_),
    .B(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4226_ (.A1(_1533_),
    .A2(_1536_),
    .A3(_1539_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4227_ (.A1(_1531_),
    .A2(_1540_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4228_ (.I(_1536_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4229_ (.I(_1539_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4230_ (.A1(_1541_),
    .A2(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4231_ (.A1(_1541_),
    .A2(_1542_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4232_ (.A1(_1533_),
    .A2(_1543_),
    .B(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4233_ (.A1(\minimax.pc_fetch[8] ),
    .A2(_1505_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4234_ (.A1(\minimax.pc_execute[8] ),
    .A2(_1504_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4235_ (.A1(_1457_),
    .A2(_1546_),
    .B(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4236_ (.A1(\minimax.regS_uc[8] ),
    .A2(_0178_),
    .B(_0078_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4237_ (.A1(_1650_),
    .A2(_1485_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4238_ (.A1(_2068_),
    .A2(_0665_),
    .B1(_1549_),
    .B2(_1403_),
    .C(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4239_ (.A1(_1548_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4240_ (.A1(_1545_),
    .A2(_1552_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4241_ (.A1(_1531_),
    .A2(_1553_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4242_ (.A1(_1548_),
    .A2(_1551_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4243_ (.A1(_1548_),
    .A2(_1551_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4244_ (.A1(_1527_),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4245_ (.A1(_1541_),
    .A2(_1542_),
    .B(_1556_),
    .C(_1519_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4246_ (.A1(_1541_),
    .A2(_1542_),
    .B1(_1548_),
    .B2(_1551_),
    .C(_1528_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4247_ (.A1(_1544_),
    .A2(_1555_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4248_ (.A1(_1554_),
    .A2(_1557_),
    .A3(_1558_),
    .A4(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4249_ (.A1(\minimax.regS_uc[9] ),
    .A2(_0178_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4250_ (.A1(_0124_),
    .A2(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4251_ (.A1(_0130_),
    .A2(_1484_),
    .B1(_1562_),
    .B2(_1433_),
    .C(_1742_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4252_ (.A1(_1550_),
    .A2(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4253_ (.A1(\minimax.pc_fetch[9] ),
    .A2(_1505_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4254_ (.A1(\minimax.pc_execute[9] ),
    .A2(_1457_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4255_ (.A1(_1458_),
    .A2(_1565_),
    .B(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4256_ (.A1(_1560_),
    .A2(_1564_),
    .A3(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4257_ (.A1(_1531_),
    .A2(_1568_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4258_ (.I(_1396_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4259_ (.A1(_1848_),
    .A2(_0641_),
    .B(_1763_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4260_ (.A1(net364),
    .A2(_0646_),
    .A3(_1415_),
    .A4(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4261_ (.A1(net386),
    .A2(net150),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4262_ (.A1(\minimax.dra[0] ),
    .A2(_1417_),
    .B1(_1572_),
    .B2(_1646_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4263_ (.A1(_1569_),
    .A2(_1571_),
    .B(_1573_),
    .C(_1387_),
    .ZN(\minimax.addrD_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4264_ (.A1(\minimax.dra[1] ),
    .A2(_1417_),
    .B1(_1572_),
    .B2(_1643_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4265_ (.A1(_1687_),
    .A2(_1571_),
    .B(_1574_),
    .ZN(\minimax.addrD_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4266_ (.A1(\minimax.dra[2] ),
    .A2(_1417_),
    .B1(_1572_),
    .B2(_0698_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4267_ (.A1(_2068_),
    .A2(_1571_),
    .B(_1575_),
    .ZN(\minimax.addrD_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4268_ (.A1(_0674_),
    .A2(_1814_),
    .B1(_1417_),
    .B2(\minimax.dra[3] ),
    .C(_1738_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4269_ (.A1(_0195_),
    .A2(_1416_),
    .B(_1576_),
    .ZN(\minimax.addrD_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4270_ (.I(\minimax.inst_regce ),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4271_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4272_ (.I(\minimax.inst_regce ),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4273_ (.A1(\inst_lat[0] ),
    .A2(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4274_ (.A1(_1851_),
    .A2(_1578_),
    .B(_1580_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4275_ (.I(_1577_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4276_ (.A1(_1581_),
    .A2(\inst_lat[1] ),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4277_ (.A1(_1626_),
    .A2(_1578_),
    .B(_1582_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4278_ (.A1(_1581_),
    .A2(\inst_lat[2] ),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4279_ (.A1(_1647_),
    .A2(_1578_),
    .B(_1583_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4280_ (.A1(_1581_),
    .A2(\inst_lat[3] ),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4281_ (.A1(_1658_),
    .A2(_1578_),
    .B(_1584_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(_1581_),
    .A2(\inst_lat[4] ),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4283_ (.A1(_1773_),
    .A2(_1578_),
    .B(_1585_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4284_ (.I(_1577_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4285_ (.A1(_1581_),
    .A2(\inst_lat[5] ),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4286_ (.A1(_0678_),
    .A2(_1586_),
    .B(_1587_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4287_ (.I(\minimax.inst_regce ),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4288_ (.A1(_1588_),
    .A2(\inst_lat[6] ),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4289_ (.A1(_1939_),
    .A2(_1586_),
    .B(_1589_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4290_ (.I0(_1396_),
    .I1(\inst_lat[7] ),
    .S(_1577_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4291_ (.I(_1590_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_1588_),
    .A2(\inst_lat[8] ),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_1687_),
    .A2(_1586_),
    .B(_1591_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4294_ (.A1(_1588_),
    .A2(\inst_lat[9] ),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4295_ (.A1(_2068_),
    .A2(_1586_),
    .B(_1592_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(_1588_),
    .A2(\inst_lat[10] ),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4297_ (.A1(_0195_),
    .A2(_1586_),
    .B(_1593_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_1577_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4299_ (.A1(_1588_),
    .A2(\inst_lat[11] ),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4300_ (.A1(_1848_),
    .A2(_1594_),
    .B(_1595_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4301_ (.A1(_1579_),
    .A2(\inst_lat[12] ),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4302_ (.A1(_1698_),
    .A2(_1594_),
    .B(_1596_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4303_ (.A1(_1579_),
    .A2(\inst_lat[13] ),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4304_ (.A1(_1812_),
    .A2(_1594_),
    .B(_1597_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4305_ (.A1(_1579_),
    .A2(\inst_lat[14] ),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4306_ (.A1(_1631_),
    .A2(_1594_),
    .B(_1598_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4307_ (.A1(_1579_),
    .A2(\inst_lat[15] ),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4308_ (.A1(_1769_),
    .A2(_1594_),
    .B(_1599_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4309_ (.A1(_1531_),
    .A2(\clknet_1_0__leaf_bank4.cen ),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4310_ (.I0(_0379_),
    .I1(\minimax.pc_fetch_dly[1] ),
    .S(_1984_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4311_ (.I(_1600_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4312_ (.I(_1634_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4313_ (.A1(\minimax.pc_fetch_dly[2] ),
    .A2(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4314_ (.A1(_1747_),
    .A2(_1602_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4315_ (.A1(\minimax.pc_fetch_dly[3] ),
    .A2(_1601_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4316_ (.A1(_1879_),
    .A2(_1603_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4317_ (.I0(\minimax.pc_fetch[4] ),
    .I1(\minimax.pc_fetch_dly[4] ),
    .S(_1984_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4318_ (.I(_1604_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4319_ (.A1(\minimax.pc_fetch_dly[5] ),
    .A2(_1601_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4320_ (.A1(_1962_),
    .A2(_1605_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4321_ (.A1(\minimax.pc_fetch_dly[6] ),
    .A2(_1601_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4322_ (.A1(_1983_),
    .A2(_1606_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(\minimax.pc_fetch_dly[7] ),
    .A2(_1601_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4324_ (.A1(_2036_),
    .A2(_1607_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4325_ (.A1(\minimax.pc_fetch_dly[8] ),
    .A2(_1749_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4326_ (.A1(_2067_),
    .A2(_1608_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4327_ (.I0(\minimax.pc_fetch[9] ),
    .I1(\minimax.pc_fetch_dly[9] ),
    .S(_1430_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4328_ (.I(_1609_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4329_ (.A1(_1531_),
    .A2(\clknet_1_0__leaf_bank3.cen ),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4330_ (.A1(_1877_),
    .A2(\clknet_1_0__leaf_bank2.cen ),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4331_ (.A1(_1877_),
    .A2(\clknet_1_0__leaf_bank1.cen ),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4332_ (.I0(\minimax.pc_fetch_dly[1] ),
    .I1(\minimax.pc_execute[1] ),
    .S(_1430_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(_1610_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4334_ (.I(_1640_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4335_ (.A1(\minimax.pc_fetch_dly[2] ),
    .A2(_1611_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4336_ (.A1(_1475_),
    .A2(_0023_),
    .B(_1612_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4337_ (.A1(\minimax.pc_fetch_dly[3] ),
    .A2(_1611_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4338_ (.A1(_1491_),
    .A2(_0023_),
    .B(_1613_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4339_ (.I(\minimax.pc_execute[4] ),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4340_ (.A1(\minimax.pc_fetch_dly[4] ),
    .A2(_1611_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4341_ (.A1(_1614_),
    .A2(_0023_),
    .B(_1615_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4342_ (.I0(\minimax.pc_fetch_dly[5] ),
    .I1(\minimax.pc_execute[5] ),
    .S(_1430_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4343_ (.I(_1616_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4344_ (.I(\minimax.pc_execute[6] ),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(\minimax.pc_fetch_dly[6] ),
    .A2(_1746_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4346_ (.A1(_1617_),
    .A2(_0023_),
    .B(_1618_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4347_ (.I(\minimax.pc_execute[7] ),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4348_ (.A1(\minimax.pc_fetch_dly[7] ),
    .A2(_1746_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4349_ (.A1(_1619_),
    .A2(_1611_),
    .B(_1620_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4350_ (.I0(\minimax.pc_fetch_dly[8] ),
    .I1(\minimax.pc_execute[8] ),
    .S(_1430_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4351_ (.I(_1621_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4352_ (.I(\minimax.pc_execute[9] ),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4353_ (.A1(\minimax.pc_fetch_dly[9] ),
    .A2(_1746_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4354_ (.A1(_1622_),
    .A2(_1611_),
    .B(_1623_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4355_ (.D(_0036_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4356_ (.D(_0037_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4357_ (.D(_0038_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4358_ (.D(_0039_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4359_ (.D(_0040_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.inst[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4360_ (.D(_0041_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.inst[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4361_ (.D(_0042_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.inst[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4362_ (.D(_0043_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.inst[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4363_ (.D(_0044_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.inst[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4364_ (.D(_0045_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.inst[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4365_ (.D(_0046_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.inst[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4366_ (.D(_0047_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4367_ (.D(_0048_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4368_ (.D(_0049_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.inst[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4369_ (.D(_0050_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4370_ (.D(_0051_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.inst[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4371_ (.D(_0018_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.dra[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4372_ (.D(_0019_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.dra[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4373_ (.D(_0020_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.dra[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4374_ (.D(_0021_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.dra[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4375_ (.D(_0022_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.dra[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4376_ (.D(\minimax.op16_lw ),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.dly16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4377_ (.D(\minimax.op16_lwsp ),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.dly16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4378_ (.D(\minimax.op16_slli_setrd ),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.dly16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4379_ (.D(\minimax.op16_slli_setrs ),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.dly16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4380_ (.D(_0023_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.inst_regce ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4381_ (.D(_0025_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4382_ (.D(_0026_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4383_ (.D(_0027_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.pc_fetch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4384_ (.D(_0028_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.pc_fetch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4385_ (.D(_0029_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.pc_fetch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4386_ (.D(_0030_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.pc_fetch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4387_ (.D(_0031_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4388_ (.D(_0032_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.pc_fetch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4389_ (.D(_0033_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _4390_ (.D(_0052_),
    .CLKN(clknet_3_6_0_wb_clk_i),
    .Q(\bank4.was_en ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4391_ (.D(_0053_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4392_ (.D(_0054_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4393_ (.D(_0055_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4394_ (.D(_0056_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4395_ (.D(_0057_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4396_ (.D(_0058_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4397_ (.D(_0059_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4398_ (.D(_0060_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4399_ (.D(_0061_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_fetch_dly[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _4400_ (.D(_0016_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.bubble1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _4401_ (.D(_0017_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\minimax.bubble2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4402_ (.D(_0024_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\minimax.microcode ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _4403_ (.D(_0062_),
    .CLKN(clknet_3_6_0_wb_clk_i),
    .Q(\bank3.was_en ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _4404_ (.D(_0063_),
    .CLKN(clknet_3_4_0_wb_clk_i),
    .Q(\bank2.was_en ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _4405_ (.D(_0064_),
    .CLKN(clknet_3_1_0_wb_clk_i),
    .Q(\bank1.was_en ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4406_ (.D(_0000_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4407_ (.D(_0007_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4408_ (.D(_0008_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4409_ (.D(_0009_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4410_ (.D(_0010_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4411_ (.D(_0011_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\inst_lat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4412_ (.D(_0012_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\inst_lat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4413_ (.D(_0013_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\inst_lat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4414_ (.D(_0014_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\inst_lat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4415_ (.D(_0015_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\inst_lat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4416_ (.D(_0001_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\inst_lat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4417_ (.D(_0002_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\inst_lat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4418_ (.D(_0003_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4419_ (.D(_0004_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\inst_lat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4420_ (.D(_0005_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4421_ (.D(_0006_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\inst_lat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4422_ (.D(_0065_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_execute[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4423_ (.D(_0066_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\minimax.pc_execute[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4424_ (.D(_0067_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.pc_execute[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4425_ (.D(_0068_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\minimax.pc_execute[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4426_ (.D(_0069_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.pc_execute[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4427_ (.D(_0070_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\minimax.pc_execute[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4428_ (.D(_0071_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_execute[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4429_ (.D(_0072_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_execute[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _4430_ (.D(_0073_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\minimax.pc_execute[9] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_16 (.I(clknet_3_0_0_wb_clk_i),
    .ZN(net359));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_15 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net358));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_14 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net357));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_13 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net356));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_12 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net355));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_11 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net354));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_10 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net353));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_9 (.I(clknet_3_2_0_wb_clk_i),
    .ZN(net352));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_8 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net351));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_7 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net350));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_6 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net349));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_5 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_4 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net347));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_3 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net346));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_2 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net345));
 gf180mcu_fd_sc_mcu7t5v0__tieh \minimax.regfile_execution_340  (.Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__tieh \minimax.regfile_execution_341  (.Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__tieh \minimax.regfile_microcode_342  (.Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__tieh \minimax.regfile_microcode_343  (.Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3255__1 (.I(clknet_3_7_0_wb_clk_i),
    .ZN(net344));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer22 (.I(net384),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer21 (.I(_1683_),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer20 (.I(_1679_),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer19 (.I(_1827_),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer18 (.I(net382),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer17 (.I(_1709_),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer16 (.I(_1770_),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer15 (.I(_1697_),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer14 (.I(_1827_),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer13 (.I(_1672_),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer12 (.I(net381),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_1827_),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer10 (.I(_0335_),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer9 (.I(_1671_),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer8 (.I(net375),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer7 (.I(net369),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer6 (.I(_1688_),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer5 (.I(net367),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer4 (.I(_1680_),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer3 (.I(net365),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer2 (.I(_1784_),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer1 (.I(_1701_),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_1__f_bank1.cen  (.I(\clknet_0_bank1.cen ),
    .Z(\clknet_1_1__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_0__f_bank1.cen  (.I(\clknet_0_bank1.cen ),
    .Z(\clknet_1_0__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_bank1.cen  (.I(\bank1.cen ),
    .Z(\clknet_0_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_1__f_bank2.cen  (.I(\clknet_0_bank2.cen ),
    .Z(\clknet_1_1__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_0__f_bank2.cen  (.I(\clknet_0_bank2.cen ),
    .Z(\clknet_1_0__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_bank2.cen  (.I(\bank2.cen ),
    .Z(\clknet_0_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_1__f_bank3.cen  (.I(\clknet_0_bank3.cen ),
    .Z(\clknet_1_1__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_0__f_bank3.cen  (.I(\clknet_0_bank3.cen ),
    .Z(\clknet_1_0__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_bank3.cen  (.I(\bank3.cen ),
    .Z(\clknet_0_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_1__f_bank4.cen  (.I(\clknet_0_bank4.cen ),
    .Z(\clknet_1_1__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_1_0__f_bank4.cen  (.I(\clknet_0_bank4.cen ),
    .Z(\clknet_1_0__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_bank4.cen  (.I(\bank4.cen ),
    .Z(\clknet_0_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_1_1_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_1_0_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_1_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_1_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_20 (.I(clknet_3_6_0_wb_clk_i),
    .ZN(net363));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_19 (.I(clknet_3_6_0_wb_clk_i),
    .ZN(net362));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_18 (.I(clknet_3_5_0_wb_clk_i),
    .ZN(net361));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_295 (.ZN(net295));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_296 (.ZN(net296));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_297 (.ZN(net297));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_331 (.ZN(net331));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_332 (.ZN(net332));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_333 (.ZN(net333));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_334 (.ZN(net334));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_335 (.ZN(net335));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_336 (.ZN(net336));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_337 (.ZN(net337));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_338 (.ZN(net338));
 gf180mcu_fd_sc_mcu7t5v0__tiel mimi_339 (.ZN(net339));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 net299_17 (.I(clknet_3_0_0_wb_clk_i),
    .ZN(net360));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4670_ (.I(net153),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4671_ (.I(net153),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4672_ (.I(net153),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4673_ (.I(net153),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4674_ (.I(net153),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4675_ (.I(net154),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4676_ (.I(net154),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4677_ (.I(net154),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(net154),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(net154),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4680_ (.I(net156),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4681_ (.I(net156),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4682_ (.I(net156),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4683_ (.I(net156),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4684_ (.I(net156),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4685_ (.I(net157),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4686_ (.I(net157),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4687_ (.I(net157),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(net161),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(net161),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(net161),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(net161),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4692_ (.I(net161),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4693_ (.I(net162),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4694_ (.I(net162),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4695_ (.I(net162),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4696_ (.I(net162),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4697_ (.I(net166),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4698_ (.I(net166),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4699_ (.I(net166),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4700_ (.I(net166),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4701_ (.I(net164),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4702_ (.I(net164),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4703_ (.I(net164),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4704_ (.I(net164),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4705_ (.I(net164),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4706_ (.I(net165),
    .Z(net63));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank1.ram1  (.CEN(\clknet_1_0__leaf_bank1.cen ),
    .CLK(net359),
    .GWEN(net148),
    .A({net118,
    net123,
    net103,
    net108,
    net133,
    net113,
    net128,
    net138,
    net143}),
    .D({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8}),
    .Q({_NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16}),
    .WEN({_NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank1.ram2  (.CEN(\clknet_1_0__leaf_bank1.cen ),
    .CLK(net358),
    .GWEN(net148),
    .A({net118,
    net123,
    net103,
    net108,
    net133,
    net113,
    net128,
    net138,
    net143}),
    .D({_NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .Q({_NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40}),
    .WEN({_NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank1.ram3  (.CEN(\clknet_1_1__leaf_bank1.cen ),
    .CLK(net357),
    .GWEN(net149),
    .A({net119,
    net124,
    net104,
    net109,
    net134,
    net114,
    net129,
    net139,
    net144}),
    .D({_NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56}),
    .Q({_NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .WEN({_NC65,
    _NC66,
    _NC67,
    _NC68,
    _NC69,
    _NC70,
    _NC71,
    _NC72}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank1.ram4  (.CEN(\clknet_1_1__leaf_bank1.cen ),
    .CLK(net356),
    .GWEN(net149),
    .A({net119,
    net124,
    net104,
    net109,
    net134,
    net114,
    net129,
    net139,
    net144}),
    .D({_NC73,
    _NC74,
    _NC75,
    _NC76,
    _NC77,
    _NC78,
    _NC79,
    _NC80}),
    .Q({_NC81,
    _NC82,
    _NC83,
    _NC84,
    _NC85,
    _NC86,
    _NC87,
    _NC88}),
    .WEN({_NC89,
    _NC90,
    _NC91,
    _NC92,
    _NC93,
    _NC94,
    _NC95,
    _NC96}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank2.ram1  (.CEN(\clknet_1_0__leaf_bank2.cen ),
    .CLK(net355),
    .GWEN(net148),
    .A({net118,
    net123,
    net103,
    net108,
    net133,
    net113,
    net128,
    net138,
    net143}),
    .D({_NC97,
    _NC98,
    _NC99,
    _NC100,
    _NC101,
    _NC102,
    _NC103,
    _NC104}),
    .Q({_NC105,
    _NC106,
    _NC107,
    _NC108,
    _NC109,
    _NC110,
    _NC111,
    _NC112}),
    .WEN({_NC113,
    _NC114,
    _NC115,
    _NC116,
    _NC117,
    _NC118,
    _NC119,
    _NC120}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank2.ram2  (.CEN(\clknet_1_0__leaf_bank2.cen ),
    .CLK(net354),
    .GWEN(net148),
    .A({net118,
    net123,
    net103,
    net108,
    net133,
    net113,
    net128,
    net138,
    net143}),
    .D({_NC121,
    _NC122,
    _NC123,
    _NC124,
    _NC125,
    _NC126,
    _NC127,
    _NC128}),
    .Q({_NC129,
    _NC130,
    _NC131,
    _NC132,
    _NC133,
    _NC134,
    _NC135,
    _NC136}),
    .WEN({_NC137,
    _NC138,
    _NC139,
    _NC140,
    _NC141,
    _NC142,
    _NC143,
    _NC144}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank2.ram3  (.CEN(\clknet_1_1__leaf_bank2.cen ),
    .CLK(net353),
    .GWEN(net149),
    .A({net119,
    net124,
    net104,
    net109,
    net134,
    net114,
    net129,
    net139,
    net144}),
    .D({_NC145,
    _NC146,
    _NC147,
    _NC148,
    _NC149,
    _NC150,
    _NC151,
    _NC152}),
    .Q({_NC153,
    _NC154,
    _NC155,
    _NC156,
    _NC157,
    _NC158,
    _NC159,
    _NC160}),
    .WEN({_NC161,
    _NC162,
    _NC163,
    _NC164,
    _NC165,
    _NC166,
    _NC167,
    _NC168}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank2.ram4  (.CEN(\clknet_1_1__leaf_bank2.cen ),
    .CLK(net352),
    .GWEN(net148),
    .A({net118,
    net123,
    net103,
    net108,
    net133,
    net113,
    net128,
    net138,
    net143}),
    .D({_NC169,
    _NC170,
    _NC171,
    _NC172,
    _NC173,
    _NC174,
    _NC175,
    _NC176}),
    .Q({_NC177,
    _NC178,
    _NC179,
    _NC180,
    _NC181,
    _NC182,
    _NC183,
    _NC184}),
    .WEN({_NC185,
    _NC186,
    _NC187,
    _NC188,
    _NC189,
    _NC190,
    _NC191,
    _NC192}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank3.ram1  (.CEN(\clknet_1_0__leaf_bank3.cen ),
    .CLK(net351),
    .GWEN(net150),
    .A({net120,
    net125,
    net105,
    net110,
    net135,
    net115,
    net130,
    net140,
    net145}),
    .D({_NC193,
    _NC194,
    _NC195,
    _NC196,
    _NC197,
    _NC198,
    _NC199,
    _NC200}),
    .Q({_NC201,
    _NC202,
    _NC203,
    _NC204,
    _NC205,
    _NC206,
    _NC207,
    _NC208}),
    .WEN({_NC209,
    _NC210,
    _NC211,
    _NC212,
    _NC213,
    _NC214,
    _NC215,
    _NC216}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank3.ram2  (.CEN(\clknet_1_0__leaf_bank3.cen ),
    .CLK(net350),
    .GWEN(net150),
    .A({net120,
    net125,
    net105,
    net110,
    net135,
    net115,
    net130,
    net140,
    net145}),
    .D({_NC217,
    _NC218,
    _NC219,
    _NC220,
    _NC221,
    _NC222,
    _NC223,
    _NC224}),
    .Q({_NC225,
    _NC226,
    _NC227,
    _NC228,
    _NC229,
    _NC230,
    _NC231,
    _NC232}),
    .WEN({_NC233,
    _NC234,
    _NC235,
    _NC236,
    _NC237,
    _NC238,
    _NC239,
    _NC240}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank3.ram3  (.CEN(\clknet_1_1__leaf_bank3.cen ),
    .CLK(net349),
    .GWEN(net151),
    .A({net121,
    net126,
    net106,
    net111,
    net136,
    net116,
    net131,
    net141,
    net146}),
    .D({_NC241,
    _NC242,
    _NC243,
    _NC244,
    _NC245,
    _NC246,
    _NC247,
    _NC248}),
    .Q({_NC249,
    _NC250,
    _NC251,
    _NC252,
    _NC253,
    _NC254,
    _NC255,
    _NC256}),
    .WEN({_NC257,
    _NC258,
    _NC259,
    _NC260,
    _NC261,
    _NC262,
    _NC263,
    _NC264}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank3.ram4  (.CEN(\clknet_1_1__leaf_bank3.cen ),
    .CLK(net348),
    .GWEN(net151),
    .A({net121,
    net126,
    net106,
    net111,
    net136,
    net116,
    net131,
    net141,
    net146}),
    .D({_NC265,
    _NC266,
    _NC267,
    _NC268,
    _NC269,
    _NC270,
    _NC271,
    _NC272}),
    .Q({_NC273,
    _NC274,
    _NC275,
    _NC276,
    _NC277,
    _NC278,
    _NC279,
    _NC280}),
    .WEN({_NC281,
    _NC282,
    _NC283,
    _NC284,
    _NC285,
    _NC286,
    _NC287,
    _NC288}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank4.ram1  (.CEN(\clknet_1_0__leaf_bank4.cen ),
    .CLK(net347),
    .GWEN(net150),
    .A({net120,
    net125,
    net105,
    net110,
    net135,
    net115,
    net130,
    net140,
    net145}),
    .D({_NC289,
    _NC290,
    _NC291,
    _NC292,
    _NC293,
    _NC294,
    _NC295,
    _NC296}),
    .Q({_NC297,
    _NC298,
    _NC299,
    _NC300,
    _NC301,
    _NC302,
    _NC303,
    _NC304}),
    .WEN({_NC305,
    _NC306,
    _NC307,
    _NC308,
    _NC309,
    _NC310,
    _NC311,
    _NC312}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank4.ram2  (.CEN(\clknet_1_0__leaf_bank4.cen ),
    .CLK(net346),
    .GWEN(net150),
    .A({net120,
    net125,
    net105,
    net110,
    net135,
    net115,
    net130,
    net140,
    net145}),
    .D({_NC313,
    _NC314,
    _NC315,
    _NC316,
    _NC317,
    _NC318,
    _NC319,
    _NC320}),
    .Q({_NC321,
    _NC322,
    _NC323,
    _NC324,
    _NC325,
    _NC326,
    _NC327,
    _NC328}),
    .WEN({_NC329,
    _NC330,
    _NC331,
    _NC332,
    _NC333,
    _NC334,
    _NC335,
    _NC336}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank4.ram3  (.CEN(\clknet_1_1__leaf_bank4.cen ),
    .CLK(net345),
    .GWEN(net151),
    .A({net121,
    net126,
    net106,
    net111,
    net136,
    net116,
    net131,
    net141,
    net146}),
    .D({_NC337,
    _NC338,
    _NC339,
    _NC340,
    _NC341,
    _NC342,
    _NC343,
    _NC344}),
    .Q({_NC345,
    _NC346,
    _NC347,
    _NC348,
    _NC349,
    _NC350,
    _NC351,
    _NC352}),
    .WEN({_NC353,
    _NC354,
    _NC355,
    _NC356,
    _NC357,
    _NC358,
    _NC359,
    _NC360}));
 gf180mcu_fd_ip_sram__sram512x8m8wm1 \bank4.ram4  (.CEN(\clknet_1_1__leaf_bank4.cen ),
    .CLK(net344),
    .GWEN(net151),
    .A({net120,
    net125,
    net105,
    net110,
    net135,
    net115,
    net130,
    net140,
    net145}),
    .D({_NC361,
    _NC362,
    _NC363,
    _NC364,
    _NC365,
    _NC366,
    _NC367,
    _NC368}),
    .Q({_NC369,
    _NC370,
    _NC371,
    _NC372,
    _NC373,
    _NC374,
    _NC375,
    _NC376}),
    .WEN({_NC377,
    _NC378,
    _NC379,
    _NC380,
    _NC381,
    _NC382,
    _NC383,
    _NC384}));
 RAM32_1RW1R \minimax.regfile_execution  (.CLK(clknet_3_4_0_wb_clk_i),
    .EN0(net340),
    .EN1(net341),
    .A0({\minimax.addrD_port[4] ,
    \minimax.addrD_port[3] ,
    \minimax.addrD_port[2] ,
    \minimax.addrD_port[1] ,
    \minimax.addrD_port[0] }),
    .A1({\minimax.addrS_port[4] ,
    \minimax.addrS_port[3] ,
    \minimax.addrS_port[2] ,
    \minimax.addrS_port[1] ,
    \minimax.addrS_port[0] }),
    .Di0({\minimax.aluX[31] ,
    \minimax.aluX[30] ,
    \minimax.aluX[29] ,
    \minimax.aluX[28] ,
    \minimax.aluX[27] ,
    \minimax.aluX[26] ,
    \minimax.aluX[25] ,
    \minimax.aluX[24] ,
    \minimax.aluX[23] ,
    \minimax.aluX[22] ,
    \minimax.aluX[21] ,
    \minimax.aluX[20] ,
    \minimax.aluX[19] ,
    \minimax.aluX[18] ,
    \minimax.aluX[17] ,
    \minimax.aluX[16] ,
    \minimax.aluX[15] ,
    \minimax.aluX[14] ,
    \minimax.aluX[13] ,
    \minimax.aluX[12] ,
    \minimax.aluX[11] ,
    \minimax.aluX[10] ,
    \minimax.aluX[9] ,
    \minimax.aluX[8] ,
    \minimax.aluX[7] ,
    \minimax.aluX[6] ,
    \minimax.aluX[5] ,
    \minimax.aluX[4] ,
    \minimax.aluX[3] ,
    \minimax.aluX[2] ,
    \minimax.aluX[1] ,
    \minimax.aluX[0] }),
    .Do0({\minimax.regD_ex[31] ,
    \minimax.regD_ex[30] ,
    \minimax.regD_ex[29] ,
    \minimax.regD_ex[28] ,
    \minimax.regD_ex[27] ,
    \minimax.regD_ex[26] ,
    \minimax.regD_ex[25] ,
    \minimax.regD_ex[24] ,
    \minimax.regD_ex[23] ,
    \minimax.regD_ex[22] ,
    \minimax.regD_ex[21] ,
    \minimax.regD_ex[20] ,
    \minimax.regD_ex[19] ,
    \minimax.regD_ex[18] ,
    \minimax.regD_ex[17] ,
    \minimax.regD_ex[16] ,
    \minimax.regD_ex[15] ,
    \minimax.regD_ex[14] ,
    \minimax.regD_ex[13] ,
    \minimax.regD_ex[12] ,
    \minimax.regD_ex[11] ,
    \minimax.regD_ex[10] ,
    \minimax.regD_ex[9] ,
    \minimax.regD_ex[8] ,
    \minimax.regD_ex[7] ,
    \minimax.regD_ex[6] ,
    \minimax.regD_ex[5] ,
    \minimax.regD_ex[4] ,
    \minimax.regD_ex[3] ,
    \minimax.regD_ex[2] ,
    \minimax.regD_ex[1] ,
    \minimax.regD_ex[0] }),
    .Do1({\minimax.regS_ex[31] ,
    \minimax.regS_ex[30] ,
    \minimax.regS_ex[29] ,
    \minimax.regS_ex[28] ,
    \minimax.regS_ex[27] ,
    \minimax.regS_ex[26] ,
    \minimax.regS_ex[25] ,
    \minimax.regS_ex[24] ,
    \minimax.regS_ex[23] ,
    \minimax.regS_ex[22] ,
    \minimax.regS_ex[21] ,
    \minimax.regS_ex[20] ,
    \minimax.regS_ex[19] ,
    \minimax.regS_ex[18] ,
    \minimax.regS_ex[17] ,
    \minimax.regS_ex[16] ,
    \minimax.regS_ex[15] ,
    \minimax.regS_ex[14] ,
    \minimax.regS_ex[13] ,
    \minimax.regS_ex[12] ,
    \minimax.regS_ex[11] ,
    \minimax.regS_ex[10] ,
    \minimax.regS_ex[9] ,
    \minimax.regS_ex[8] ,
    \minimax.regS_ex[7] ,
    \minimax.regS_ex[6] ,
    \minimax.regS_ex[5] ,
    \minimax.regS_ex[4] ,
    \minimax.regS_ex[3] ,
    \minimax.regS_ex[2] ,
    \minimax.regS_ex[1] ,
    \minimax.regS_ex[0] }),
    .WE0({_0034_,
    _0034_,
    _0034_,
    _0034_}));
 RAM32_1RW1R \minimax.regfile_microcode  (.CLK(clknet_3_7_0_wb_clk_i),
    .EN0(net342),
    .EN1(net343),
    .A0({\minimax.addrD_port[4] ,
    \minimax.addrD_port[3] ,
    \minimax.addrD_port[2] ,
    \minimax.addrD_port[1] ,
    \minimax.addrD_port[0] }),
    .A1({\minimax.addrS_port[4] ,
    \minimax.addrS_port[3] ,
    \minimax.addrS_port[2] ,
    \minimax.addrS_port[1] ,
    \minimax.addrS_port[0] }),
    .Di0({\minimax.aluX[31] ,
    \minimax.aluX[30] ,
    \minimax.aluX[29] ,
    \minimax.aluX[28] ,
    \minimax.aluX[27] ,
    \minimax.aluX[26] ,
    \minimax.aluX[25] ,
    \minimax.aluX[24] ,
    \minimax.aluX[23] ,
    \minimax.aluX[22] ,
    \minimax.aluX[21] ,
    \minimax.aluX[20] ,
    \minimax.aluX[19] ,
    \minimax.aluX[18] ,
    \minimax.aluX[17] ,
    \minimax.aluX[16] ,
    \minimax.aluX[15] ,
    \minimax.aluX[14] ,
    \minimax.aluX[13] ,
    \minimax.aluX[12] ,
    \minimax.aluX[11] ,
    \minimax.aluX[10] ,
    \minimax.aluX[9] ,
    \minimax.aluX[8] ,
    \minimax.aluX[7] ,
    \minimax.aluX[6] ,
    \minimax.aluX[5] ,
    \minimax.aluX[4] ,
    \minimax.aluX[3] ,
    \minimax.aluX[2] ,
    \minimax.aluX[1] ,
    \minimax.aluX[0] }),
    .Do0({\minimax.regD_uc[31] ,
    \minimax.regD_uc[30] ,
    \minimax.regD_uc[29] ,
    \minimax.regD_uc[28] ,
    \minimax.regD_uc[27] ,
    \minimax.regD_uc[26] ,
    \minimax.regD_uc[25] ,
    \minimax.regD_uc[24] ,
    \minimax.regD_uc[23] ,
    \minimax.regD_uc[22] ,
    \minimax.regD_uc[21] ,
    \minimax.regD_uc[20] ,
    \minimax.regD_uc[19] ,
    \minimax.regD_uc[18] ,
    \minimax.regD_uc[17] ,
    \minimax.regD_uc[16] ,
    \minimax.regD_uc[15] ,
    \minimax.regD_uc[14] ,
    \minimax.regD_uc[13] ,
    \minimax.regD_uc[12] ,
    \minimax.regD_uc[11] ,
    \minimax.regD_uc[10] ,
    \minimax.regD_uc[9] ,
    \minimax.regD_uc[8] ,
    \minimax.regD_uc[7] ,
    \minimax.regD_uc[6] ,
    \minimax.regD_uc[5] ,
    \minimax.regD_uc[4] ,
    \minimax.regD_uc[3] ,
    \minimax.regD_uc[2] ,
    \minimax.regD_uc[1] ,
    \minimax.regD_uc[0] }),
    .Do1({\minimax.regS_uc[31] ,
    \minimax.regS_uc[30] ,
    \minimax.regS_uc[29] ,
    \minimax.regS_uc[28] ,
    \minimax.regS_uc[27] ,
    \minimax.regS_uc[26] ,
    \minimax.regS_uc[25] ,
    \minimax.regS_uc[24] ,
    \minimax.regS_uc[23] ,
    \minimax.regS_uc[22] ,
    \minimax.regS_uc[21] ,
    \minimax.regS_uc[20] ,
    \minimax.regS_uc[19] ,
    \minimax.regS_uc[18] ,
    \minimax.regS_uc[17] ,
    \minimax.regS_uc[16] ,
    \minimax.regS_uc[15] ,
    \minimax.regS_uc[14] ,
    \minimax.regS_uc[13] ,
    \minimax.regS_uc[12] ,
    \minimax.regS_uc[11] ,
    \minimax.regS_uc[10] ,
    \minimax.regS_uc[9] ,
    \minimax.regS_uc[8] ,
    \minimax.regS_uc[7] ,
    \minimax.regS_uc[6] ,
    \minimax.regS_uc[5] ,
    \minimax.regS_uc[4] ,
    \minimax.regS_uc[3] ,
    \minimax.regS_uc[2] ,
    \minimax.regS_uc[1] ,
    \minimax.regS_uc[0] }),
    .WE0({_0035_,
    _0035_,
    _0035_,
    _0035_}));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_15999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_16773 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1 (.I(wb_rst_i),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input2 (.I(wbs_dat_i[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input3 (.I(wbs_dat_i[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input4 (.I(wbs_dat_i[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input5 (.I(wbs_dat_i[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input6 (.I(wbs_dat_i[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input7 (.I(wbs_dat_i[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input8 (.I(wbs_dat_i[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input9 (.I(wbs_dat_i[16]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input10 (.I(wbs_dat_i[17]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input11 (.I(wbs_dat_i[18]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input12 (.I(wbs_dat_i[19]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input13 (.I(wbs_dat_i[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input14 (.I(wbs_dat_i[20]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input15 (.I(wbs_dat_i[21]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input16 (.I(wbs_dat_i[22]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input17 (.I(wbs_dat_i[23]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input18 (.I(wbs_dat_i[24]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input19 (.I(wbs_dat_i[25]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input20 (.I(wbs_dat_i[26]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input21 (.I(wbs_dat_i[27]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 input22 (.I(wbs_dat_i[28]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input23 (.I(wbs_dat_i[29]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input24 (.I(wbs_dat_i[2]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input25 (.I(wbs_dat_i[30]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input26 (.I(wbs_dat_i[31]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input27 (.I(wbs_dat_i[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input28 (.I(wbs_dat_i[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(wbs_dat_i[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(wbs_dat_i[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(wbs_dat_i[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(wbs_dat_i[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(wbs_dat_i[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(io_oeb[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(io_oeb[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(io_oeb[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(io_oeb[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(io_oeb[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(io_oeb[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(io_oeb[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(io_oeb[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(io_oeb[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(io_oeb[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(io_oeb[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(io_oeb[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(io_oeb[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(io_oeb[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(io_oeb[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(io_oeb[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(io_oeb[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output80 (.I(net80),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output81 (.I(net81),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output82 (.I(net82),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output84 (.I(net84),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output85 (.I(net85),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output86 (.I(net86),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output87 (.I(net87),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output88 (.I(net88),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output89 (.I(net89),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output90 (.I(net90),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output91 (.I(net91),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output92 (.I(net92),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output93 (.I(net93),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output94 (.I(net94),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output95 (.I(net95),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output96 (.I(net96),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output97 (.I(net97),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output98 (.I(net98),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output99 (.I(net99),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output100 (.I(net100),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output101 (.I(net101),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output102 (.I(net102),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout103 (.I(net107),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout104 (.I(net107),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout105 (.I(net107),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout107 (.I(\bank1.addr[6] ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout108 (.I(net112),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout109 (.I(net112),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout110 (.I(net112),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout112 (.I(\bank1.addr[5] ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout113 (.I(net117),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout114 (.I(net117),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout115 (.I(net117),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout117 (.I(\bank1.addr[3] ),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout118 (.I(net122),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout119 (.I(net122),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout120 (.I(net122),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout122 (.I(\bank1.addr[8] ),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout123 (.I(net127),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout124 (.I(net127),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout125 (.I(net127),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout127 (.I(\bank1.addr[7] ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout128 (.I(net132),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout129 (.I(net132),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout130 (.I(net132),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout132 (.I(\bank1.addr[2] ),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout133 (.I(net137),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout134 (.I(net137),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout135 (.I(net137),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout137 (.I(\bank1.addr[4] ),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout138 (.I(net142),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout139 (.I(net142),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout140 (.I(net142),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout142 (.I(\bank1.addr[1] ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout143 (.I(net147),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout144 (.I(net147),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout145 (.I(net147),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout146 (.I(net147),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout147 (.I(\bank1.addr[0] ),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout148 (.I(net152),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 fanout149 (.I(net152),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_16 fanout150 (.I(net152),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 fanout151 (.I(net152),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 fanout152 (.I(\bank1.wen_mask[0] ),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout153 (.I(net155),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout154 (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout155 (.I(net159),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout156 (.I(net158),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout157 (.I(net158),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout158 (.I(net159),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout159 (.I(net160),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 fanout160 (.I(net168),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout161 (.I(net163),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout162 (.I(net163),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout163 (.I(net167),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout164 (.I(net165),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout165 (.I(net166),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout166 (.I(net167),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout167 (.I(net168),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 fanout168 (.I(net1),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer23 (.I(_1825_),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer24 (.I(net386),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer25 (.I(_2013_),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer26 (.I(_1751_),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer27 (.I(_1828_),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer28 (.I(_1678_),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer29 (.I(net391),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer30 (.I(net392),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer31 (.I(_1714_),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer32 (.I(net394),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer33 (.I(_0349_),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer34 (.I(_1718_),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer35 (.I(_1663_),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer36 (.I(net398),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer37 (.I(_1970_),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer38 (.I(_1713_),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer39 (.I(_0336_),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer40 (.I(_0305_),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer41 (.I(_1828_),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer42 (.I(_1942_),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 rebuffer43 (.I(_1670_),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer44 (.I(net406),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer45 (.I(_1699_),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer46 (.I(_0129_),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer47 (.I(\minimax.inst[10] ),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer48 (.I(net410),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__D (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__D (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__D (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__D (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__D (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__D (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__D (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__D (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__D (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__D (.I(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__D (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__D (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_WE0[3]  (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_WE0[2]  (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_WE0[1]  (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_WE0[0]  (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_WE0[3]  (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_WE0[2]  (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_WE0[1]  (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_WE0[0]  (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__D (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__D (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__D (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__I (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__B (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__B1 (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__I (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__S (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__S (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__S (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__S (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A3 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A3 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A3 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A3 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A4 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__B (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A2 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A3 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__I (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__B (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__I (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__B2 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A2 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__C (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A1 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A3 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A3 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B2 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__I (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__B2 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__B (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__B (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__B (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A2 (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A3 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A1 (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__I (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A3 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A3 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B3 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__I (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__I (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A3 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A1 (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A3 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__C (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A2 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__B (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__C (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer46_I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A3 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__B2 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__B2 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__B2 (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__B (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__B (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A2 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A2 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__B (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A2 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A3 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__B (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__A1 (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A3 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__I (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__B1 (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A1 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__B2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A2 (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A2 (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__I (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A2 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__C (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__C (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__I (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A2 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__B (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__B (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__C (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__B2 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__I (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__B (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__B2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__B2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__I (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__C (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A2 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__B (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__B2 (.I(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A2 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__I (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__S (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__S (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__S (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__I (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__I (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A2 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A3 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__B (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A4 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__A1 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A1 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__I (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__B (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__S (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__S (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__I (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__B2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__B2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__I (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__B2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A2 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__A2 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__I (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A4 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A2 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__B1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__I (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__B (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__B2 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A2 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__B (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__I (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__I (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__B (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__B (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__B (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__B (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__I (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__I (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__B2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A1 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__I0 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__I1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__I (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A2 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A3 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__I (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A3 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__A2 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__B (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A3 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A4 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A3 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A3 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A3 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A3 (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A3 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A1 (.I(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3310__I (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3306__I (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__B2 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__A1 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A2 (.I(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A3 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A3 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A3 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A4 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A3 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A3 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A4 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A2 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__B (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__I (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__I (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__I (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A4 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A3 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A2 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A2 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A3 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__B2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A2 (.I(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A3 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A3 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A3 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A3 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__A3 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2861__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__S (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__I (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__I (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__B (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__A2 (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__B (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__I (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__I (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A3 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A4 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A2 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A3 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A4 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__B (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__B1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A3 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A3 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A4 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__A3 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__B (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__C (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__B (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3354__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__B (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__C (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2867__B (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__A4 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A3 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__B2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B2 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__C (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__A1 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A3 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__B (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__B (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__I (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__B (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__C (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer40_I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A3 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A3 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__B (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A4 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A3 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__B (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2873__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__B2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__B1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A3 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A3 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__C (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__B (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__B (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer10_I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer39_I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A3 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2895__A2 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__I (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A3 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A3 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3113__S (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__B (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__B (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3001__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__B (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__B (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2941__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__B (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__B (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__B (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__B (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__B (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3013__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A3 (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__I (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I0 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__S (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__S (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__I (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__B (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__B (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__B (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__B1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3046__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__B2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__B (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__B (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__B (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__B (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__B (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3136__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3025__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__I (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A1 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__I (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__S (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__S (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__S (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__S (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__B (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__B2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__I (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__S (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__S (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__S (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__B2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__B2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__B2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__B2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__B2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__B2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3026__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3027__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__I (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__C2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__I (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3072__I (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3080__I (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__S (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__C (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__B (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__C (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A3 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3172__A3 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__A3 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A3 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A2 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__B2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__A2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3117__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__I (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__I (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A3 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__B2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__I (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__B (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__B (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__A3 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A3 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__S (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__S (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__S (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__S (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__S (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3230__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3252__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A3 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__B2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__B (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A3 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__I0 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__A2 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__B1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A3 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A3 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__B2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__B2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__S (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__C (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__B2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__B (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__A3 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A3 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__B1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__B2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3352__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__B (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A3 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__B2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A3 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__B (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A4 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3308__A2 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__C (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__B2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3312__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__I0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__I0 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3316__A3 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__A3 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__C (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__C (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__C (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__I (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__C (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3395__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__B (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__B1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A2 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__I1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A3 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__B2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__B2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__B (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__A3 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3399__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A3 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__C1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__C1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__C1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__B1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__B (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__B (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__B1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__B2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3356__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__B (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__B (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__I (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A3 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A3 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__B1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__B2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__B1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__B2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__C (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__B (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__B (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__B (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__B (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__A3 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A3 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__I1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__I1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I0 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3397__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__C (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__B1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__C (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__C (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__B1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__B2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__B2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__C (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__B2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__B2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A3 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__B1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__B2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__B (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__B (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__I0 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I0 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A3 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A3 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__C (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__B (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__C1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__B1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__B2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__B2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__B2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__C (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__B (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__B1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__B2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__B (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__B2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__B (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__C (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__B (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__S (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__S (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__S (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__B (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__B (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__B (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__B (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A3 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A3 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I0 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__A3 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A4 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__B2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__B (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__B2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A3 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__B2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__B2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__C (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__C (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__B2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__C (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__B1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__C (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A3 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A3 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__B1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A2 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A3 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__I0 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__B1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A3 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__B2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__C (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__C (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A4 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A4 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A4 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A4 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__C (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A3 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__B1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__B2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__B (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__I (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A3 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A2 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A4 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__I (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__S (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A3 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__B1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__C (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__B1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A3 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__C (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__B (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__B1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I0 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__C (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A3 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A3 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__B (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__C (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A3 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A3 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A4 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__B (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3606__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__B (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__C (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__B (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__B (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A3 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__C (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__B (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__C (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A4 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A2 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__B (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I0 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A4 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A4 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A3 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__B (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__B (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A3 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__B (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A3 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__C (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__B (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__S (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__S (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A3 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A3 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__B2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A3 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A3 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A3 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__B (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__B (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__B (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__B (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__B (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A3 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__B2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__B1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A4 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__A3 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__B2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__C (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__B (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3709__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A3 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__S (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__B (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__B1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A4 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__C (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A2 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__C (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__B (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__I1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A3 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A3 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A3 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A4 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I0 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A4 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A4 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__S (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__S (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__S (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__C (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A3 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__B (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__C (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3759__A3 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__B (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__C (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__B (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__C (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__C (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__I (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__B (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__B1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A4 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__C (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A3 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__B (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__B2 (.I(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__B (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__S (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__C (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__I0 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__I1 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A3 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A3 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I0 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A4 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A3 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A3 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A4 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A3 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__B (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__B2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__B2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A3 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__C (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__C (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A3 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__A3 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__A3 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__C (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A3 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__B1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__I (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__B (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A3 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__B2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A3 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__B1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__B1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__B (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__B (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__C (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__B (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__B (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A3 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A3 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__I (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A3 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__B1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__B (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__C (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__B (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__C (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A3 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A3 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__I (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A3 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A3 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A4 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A3 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A4 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__B (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A3 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A3 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A4 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A3 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__B1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__B (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__C (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__B (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__C (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__B (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__C (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__B1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__B2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__B2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__S (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__B (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__C (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__C (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__C (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__C (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__B2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__B (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__B (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__B1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A3 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__C (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__B (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__B1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__B1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__I0 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__I (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__B2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__C1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__C (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__B (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__B (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__B (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A3 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__I (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__B2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__B (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B (.I(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B1 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__B (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__C2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__C2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__C (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__I (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A3 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A3 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__B1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__B (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__B1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__B1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__B1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__S (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__S (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__S (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__S (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A3 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__B2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__B2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A3 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A3 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A3 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A3 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A3 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A3 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__S (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__S (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__B1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A4 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A3 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A3 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A4 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__I (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A3 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__I1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__B1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__B1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__C (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__I1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A3 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__B (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__C (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__C (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__C (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__B (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__B (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__B1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__I (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__B1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__B1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__C (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__B2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__B1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__B (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__B (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__S (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__B (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__B (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__B (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__B (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__B (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__B (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__B (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__B (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__B (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__B (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__B (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__B (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__B (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__B (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__B (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__B (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__I (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__I (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__B (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A1 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__B (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__B2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__I (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A3 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A3 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__I (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__B2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__B2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__B2 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B2 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__B (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__C (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__I (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__C (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__B (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A3 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__B (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A4 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A3 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A3 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A2 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A3 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__I (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A3 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A3 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__I (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A4 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A4 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A3 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__I (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__I (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer35_I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A3 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A3 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__B2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__I (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__I (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__I (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer43_I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A3 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer9_I (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A3 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A4 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer13_I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__B2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A3 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__A3 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__I1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A4 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__S (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__I (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__I (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer28_I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A4 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer20_I (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A3 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A3 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer4_I (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__C (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__B1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer21_I (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__C (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__I (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A3 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer6_I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A3 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__A3 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__I (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A4 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A4 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A4 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A3 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A4 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__I (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A3 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A3 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__B (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer15_I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer45_I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__B1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A3 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer1_I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__C2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__C1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A3 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A3 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer17_I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A3 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A3 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer38_I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__A3 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer31_I (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__B1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__I (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A3 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A3 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A3 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A3 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__I (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A3 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A3 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A3 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__S (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__S (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__S (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__B1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__S (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__I (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__S (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__S (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__I (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__S (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__S (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__S (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__S (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__S (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__S (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__S (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__S (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__I (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__S (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__S (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__S (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__I (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__I (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__S (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__S (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__S (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__I (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__C (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A3 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A3 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A3 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__I (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__C (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A3 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__I (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__B2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer26_I (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A4 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A2 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__B (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__I (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__I (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__B (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A3 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A3 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__I (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__B (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I0 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__I (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__B (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__B (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__A1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A3 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__I (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__I (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__I (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__B2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A4 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__I (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__B2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A3 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer16_I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A3 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A4 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__I (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__I (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__C (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A3 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__B (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A2 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__B (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__I (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A3 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__I (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__I (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__B (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__S (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__S (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__S (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__I0 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__S (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__B2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__I1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A2 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A2 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__B2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__I (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__I (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__B1 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__C1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__I (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__B2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__S (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__S (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__C (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer19_I (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer14_I (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer11_I (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer41_I (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer27_I (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A3 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A3 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__I (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A3 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__I (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__B2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__B2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__B2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__B (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__B1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__C (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__I (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A3 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__I (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A3 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__B (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__I (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A3 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A3 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__B1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__B (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__I (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__B2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__B (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A3 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A3 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__B (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A3 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A3 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A3 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__S (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__B (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A1 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__C (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A1 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__B1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A3 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A4 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__A3 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A3 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__I1 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A4 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__A1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__B1 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__B2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__B1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__B2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__B (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__B1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3425__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__B1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__I (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__I (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__I (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__B (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__B (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__B (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__I (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__B2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3358__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__I (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__B2 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A1 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__B (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__I (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__B (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3362__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A3 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__B (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__B (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__I (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__C (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__I (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A3 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__B1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__C1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__B (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__I (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A3 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A3 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__I (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A3 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A3 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A3 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A3 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__I (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__B (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A3 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A4 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A4 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A3 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3318__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__C (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__C (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer42_I (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__I (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__B (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__B2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A4 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__B (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A3 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A4 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__B (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3374__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__C (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A1 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B1 (.I(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__B (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__I (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__I (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer37_I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A3 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A3 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A3 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__I (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A3 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A4 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__C (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A3 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__B (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__B2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__I (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2528__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__S (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__S (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__I (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__A1 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__A1 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A3 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A3 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__B2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__C (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__C (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3372__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__B (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__I (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__A1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I0 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__I (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer25_I (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__B (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__C (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__B2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__I (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__S (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__C (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__I (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__B (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__C (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A4 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A4 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__I (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__I (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__B (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__B (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__B (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__B (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__S (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__S (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__S (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__S (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__I (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__I (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A3 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__B2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__B2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A3 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A3 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__B1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__B (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__I (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__B2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__B2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__B (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__B1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__B (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__B1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__I (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__I (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A1 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__I (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__A2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__A3 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A4 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__I (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A3 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__B (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__A4 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A3 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A3 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A3 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A3 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__B2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A3 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__I (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B2 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__I (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__S (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__I (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__I (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__I0 (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A2 (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A3 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A2 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__I (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__A1 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(net364));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_CEN  (.I(\clknet_1_1__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_CEN  (.I(\clknet_1_1__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A2 (.I(\clknet_1_0__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_CEN  (.I(\clknet_1_0__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_CEN  (.I(\clknet_1_0__leaf_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_1__f_bank1.cen_I  (.I(\clknet_0_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_0__f_bank1.cen_I  (.I(\clknet_0_bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_CEN  (.I(\clknet_1_1__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_CEN  (.I(\clknet_1_1__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(\clknet_1_0__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_CEN  (.I(\clknet_1_0__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_CEN  (.I(\clknet_1_0__leaf_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_1__f_bank2.cen_I  (.I(\clknet_0_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_0__f_bank2.cen_I  (.I(\clknet_0_bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_CEN  (.I(\clknet_1_1__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_CEN  (.I(\clknet_1_1__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(\clknet_1_0__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_CEN  (.I(\clknet_1_0__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_CEN  (.I(\clknet_1_0__leaf_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_1__f_bank3.cen_I  (.I(\clknet_0_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_0__f_bank3.cen_I  (.I(\clknet_0_bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_CEN  (.I(\clknet_1_1__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_CEN  (.I(\clknet_1_1__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(\clknet_1_0__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_CEN  (.I(\clknet_1_0__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_CEN  (.I(\clknet_1_0__leaf_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_1__f_bank4.cen_I  (.I(\clknet_0_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_1_0__f_bank4.cen_I  (.I(\clknet_0_bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_CLK  (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3255__1_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_2_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_3_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_4_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_5_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_6_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_7_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_8_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__CLKN (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__CLKN (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_19_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_20_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_18_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__CLKN (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_CLK  (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_9_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_10_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_11_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_12_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_13_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_14_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_15_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__CLKN (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_16_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_net299_17_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_1_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_1_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(\bank1.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(\bank1.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(\bank1.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(\bank1.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(\bank1.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(\bank1.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(\bank1.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(\bank1.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(\bank1.addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_bank1.cen_I  (.I(\bank1.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(\bank1.rdata[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A1 (.I(\bank1.rdata[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(\bank1.rdata[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A1 (.I(\bank1.rdata[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(\bank1.rdata[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(\bank1.rdata[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__A1 (.I(\bank1.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A1 (.I(\bank1.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A1 (.I(\bank1.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__A1 (.I(\bank1.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3378__A1 (.I(\bank1.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(\bank1.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(\bank1.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__A1 (.I(\bank1.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(\bank1.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__A1 (.I(\bank1.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__A1 (.I(\bank1.rdata[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__A1 (.I(\bank1.rdata[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(\bank1.wen_mask[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_bank2.cen_I  (.I(\bank2.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__A1 (.I(\bank2.was_en ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_bank3.cen_I  (.I(\bank3.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_bank4.cen_I  (.I(\bank4.cen ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(\inst_lat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(\inst_lat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(\inst_lat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(\inst_lat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(\inst_lat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(\inst_lat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(\inst_lat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(\inst_lat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(\inst_lat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(\inst_lat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(\inst_lat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A2 (.I(\inst_lat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A2 (.I(\inst_lat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__I1 (.I(\inst_lat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(\inst_lat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(\inst_lat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A0[0]  (.I(\minimax.addrD_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A0[0]  (.I(\minimax.addrD_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A0[1]  (.I(\minimax.addrD_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A0[1]  (.I(\minimax.addrD_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A0[2]  (.I(\minimax.addrD_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A0[2]  (.I(\minimax.addrD_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A0[3]  (.I(\minimax.addrD_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A0[3]  (.I(\minimax.addrD_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A0[4]  (.I(\minimax.addrD_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A0[4]  (.I(\minimax.addrD_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A1[0]  (.I(\minimax.addrS_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A1[0]  (.I(\minimax.addrS_port[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A1[1]  (.I(\minimax.addrS_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A1[1]  (.I(\minimax.addrS_port[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A1[2]  (.I(\minimax.addrS_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A1[2]  (.I(\minimax.addrS_port[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A1[3]  (.I(\minimax.addrS_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A1[3]  (.I(\minimax.addrS_port[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_A1[4]  (.I(\minimax.addrS_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_A1[4]  (.I(\minimax.addrS_port[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[0]  (.I(\minimax.aluX[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[0]  (.I(\minimax.aluX[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[10]  (.I(\minimax.aluX[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[10]  (.I(\minimax.aluX[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[11]  (.I(\minimax.aluX[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[11]  (.I(\minimax.aluX[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[12]  (.I(\minimax.aluX[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[12]  (.I(\minimax.aluX[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[13]  (.I(\minimax.aluX[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[13]  (.I(\minimax.aluX[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[14]  (.I(\minimax.aluX[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[14]  (.I(\minimax.aluX[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[15]  (.I(\minimax.aluX[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[15]  (.I(\minimax.aluX[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[16]  (.I(\minimax.aluX[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[16]  (.I(\minimax.aluX[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[17]  (.I(\minimax.aluX[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[17]  (.I(\minimax.aluX[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[18]  (.I(\minimax.aluX[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[18]  (.I(\minimax.aluX[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[19]  (.I(\minimax.aluX[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[19]  (.I(\minimax.aluX[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[1]  (.I(\minimax.aluX[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[1]  (.I(\minimax.aluX[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[20]  (.I(\minimax.aluX[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[20]  (.I(\minimax.aluX[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[21]  (.I(\minimax.aluX[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[21]  (.I(\minimax.aluX[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[22]  (.I(\minimax.aluX[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[22]  (.I(\minimax.aluX[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[23]  (.I(\minimax.aluX[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[23]  (.I(\minimax.aluX[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[24]  (.I(\minimax.aluX[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[24]  (.I(\minimax.aluX[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[25]  (.I(\minimax.aluX[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[25]  (.I(\minimax.aluX[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[26]  (.I(\minimax.aluX[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[26]  (.I(\minimax.aluX[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[27]  (.I(\minimax.aluX[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[27]  (.I(\minimax.aluX[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[28]  (.I(\minimax.aluX[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[28]  (.I(\minimax.aluX[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[29]  (.I(\minimax.aluX[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[29]  (.I(\minimax.aluX[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[2]  (.I(\minimax.aluX[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[2]  (.I(\minimax.aluX[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[30]  (.I(\minimax.aluX[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[30]  (.I(\minimax.aluX[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[31]  (.I(\minimax.aluX[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[31]  (.I(\minimax.aluX[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[3]  (.I(\minimax.aluX[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[3]  (.I(\minimax.aluX[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[4]  (.I(\minimax.aluX[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[4]  (.I(\minimax.aluX[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[5]  (.I(\minimax.aluX[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[5]  (.I(\minimax.aluX[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[6]  (.I(\minimax.aluX[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[6]  (.I(\minimax.aluX[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[7]  (.I(\minimax.aluX[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[7]  (.I(\minimax.aluX[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[8]  (.I(\minimax.aluX[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[8]  (.I(\minimax.aluX[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_microcode_Di0[9]  (.I(\minimax.aluX[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_minimax.regfile_execution_Di0[9]  (.I(\minimax.aluX[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A2 (.I(\minimax.dly16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A2 (.I(\minimax.dly16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(\minimax.dly16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(\minimax.dly16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(\minimax.dly16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(\minimax.dly16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(\minimax.dly16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A2 (.I(\minimax.dly16_slli_setrd ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__I (.I(\minimax.dly16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__I (.I(\minimax.dly16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A2 (.I(\minimax.dly16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2324__A2 (.I(\minimax.dly16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A1 (.I(\minimax.dra[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(\minimax.dra[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(\minimax.dra[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(\minimax.dra[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(\minimax.dra[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(\minimax.dra[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__B2 (.I(\minimax.dra[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(\minimax.dra[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B2 (.I(\minimax.dra[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(\minimax.dra[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__I (.I(\minimax.inst[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(\minimax.inst[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__I (.I(\minimax.inst[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(\minimax.inst[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A4 (.I(\minimax.inst[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__I (.I(\minimax.inst[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A2 (.I(\minimax.inst[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(\minimax.inst[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__I (.I(\minimax.inst[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__I (.I(\minimax.inst[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(\minimax.inst[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(\minimax.inst[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__C (.I(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__I (.I(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__A2 (.I(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__I (.I(\minimax.inst[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__I (.I(\minimax.inst[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__I (.I(\minimax.inst[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__I (.I(\minimax.inst[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(\minimax.inst[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__I (.I(\minimax.inst[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__I (.I(\minimax.inst[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(\minimax.inst[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__I (.I(\minimax.inst[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__A2 (.I(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__I (.I(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__I (.I(\minimax.inst[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__I (.I(\minimax.inst[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A2 (.I(\minimax.inst[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I (.I(\minimax.inst[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A3 (.I(\minimax.inst[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__I (.I(\minimax.inst[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__C2 (.I(\minimax.inst[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A1 (.I(\minimax.inst[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(\minimax.inst[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__I (.I(\minimax.inst[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A2 (.I(\minimax.inst[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A2 (.I(\minimax.inst[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__I (.I(\minimax.inst_regce ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(\minimax.inst_regce ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__I (.I(\minimax.inst_regce ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(\minimax.microcode ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A1 (.I(\minimax.microcode ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(\minimax.microcode ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__D (.I(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__C (.I(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(\minimax.op16_lw ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__D (.I(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(\minimax.op16_lwsp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__D (.I(\minimax.op16_slli_setrs ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I1 (.I(\minimax.pc_execute[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(\minimax.pc_execute[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(\minimax.pc_execute[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__I (.I(\minimax.pc_execute[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(\minimax.pc_execute[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__I (.I(\minimax.pc_execute[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(\minimax.pc_execute[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I1 (.I(\minimax.pc_execute[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(\minimax.pc_execute[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I1 (.I(\minimax.pc_execute[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(\minimax.pc_execute[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(\minimax.pc_fetch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(\minimax.pc_fetch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__I (.I(\minimax.pc_fetch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__I (.I(\minimax.pc_fetch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(\minimax.pc_fetch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(\minimax.pc_fetch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(\minimax.pc_fetch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(\minimax.pc_fetch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I0 (.I(\minimax.pc_fetch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(\minimax.pc_fetch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(\minimax.pc_fetch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(\minimax.pc_fetch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(\minimax.pc_fetch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(\minimax.pc_fetch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(\minimax.pc_fetch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(\minimax.pc_fetch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(\minimax.pc_fetch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(\minimax.pc_fetch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(\minimax.pc_fetch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I0 (.I(\minimax.pc_fetch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(\minimax.pc_fetch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(\minimax.pc_fetch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I0 (.I(\minimax.pc_fetch_dly[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I1 (.I(\minimax.pc_fetch_dly[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__B2 (.I(\minimax.pc_fetch_dly[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(\minimax.pc_fetch_dly[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(\minimax.pc_fetch_dly[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__B2 (.I(\minimax.pc_fetch_dly[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(\minimax.pc_fetch_dly[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(\minimax.pc_fetch_dly[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__C2 (.I(\minimax.pc_fetch_dly[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A1 (.I(\minimax.pc_fetch_dly[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I1 (.I(\minimax.pc_fetch_dly[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__C2 (.I(\minimax.pc_fetch_dly[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I0 (.I(\minimax.pc_fetch_dly[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(\minimax.pc_fetch_dly[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__C2 (.I(\minimax.pc_fetch_dly[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(\minimax.pc_fetch_dly[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(\minimax.pc_fetch_dly[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__B2 (.I(\minimax.pc_fetch_dly[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(\minimax.pc_fetch_dly[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(\minimax.pc_fetch_dly[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__B2 (.I(\minimax.pc_fetch_dly[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I0 (.I(\minimax.pc_fetch_dly[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(\minimax.pc_fetch_dly[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__B2 (.I(\minimax.pc_fetch_dly[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A1 (.I(\minimax.pc_fetch_dly[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I1 (.I(\minimax.pc_fetch_dly[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__B2 (.I(\minimax.pc_fetch_dly[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(\minimax.regD_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__I0 (.I(\minimax.regD_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I0 (.I(\minimax.regD_ex[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I0 (.I(\minimax.regD_ex[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__I0 (.I(\minimax.regD_ex[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I0 (.I(\minimax.regD_ex[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__I0 (.I(\minimax.regD_ex[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(\minimax.regD_ex[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__I0 (.I(\minimax.regD_ex[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__I0 (.I(\minimax.regD_ex[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__I0 (.I(\minimax.regD_ex[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__I0 (.I(\minimax.regD_ex[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(\minimax.regD_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A1 (.I(\minimax.regD_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(\minimax.regD_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__I0 (.I(\minimax.regD_ex[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__I0 (.I(\minimax.regD_ex[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__I0 (.I(\minimax.regD_ex[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__I0 (.I(\minimax.regD_ex[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I0 (.I(\minimax.regD_ex[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__I0 (.I(\minimax.regD_ex[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__I0 (.I(\minimax.regD_ex[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__I0 (.I(\minimax.regD_ex[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__I0 (.I(\minimax.regD_ex[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__I0 (.I(\minimax.regD_ex[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(\minimax.regD_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__I0 (.I(\minimax.regD_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__I0 (.I(\minimax.regD_ex[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__I0 (.I(\minimax.regD_ex[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__I0 (.I(\minimax.regD_ex[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__I0 (.I(\minimax.regD_ex[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__I0 (.I(\minimax.regD_ex[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A1 (.I(\minimax.regD_ex[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__I0 (.I(\minimax.regD_ex[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I0 (.I(\minimax.regD_ex[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__I0 (.I(\minimax.regD_ex[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(\minimax.regD_ex[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(\minimax.regD_ex[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I0 (.I(\minimax.regD_ex[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A1 (.I(\minimax.regD_ex[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__I0 (.I(\minimax.regD_ex[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(\minimax.regD_ex[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__I0 (.I(\minimax.regD_ex[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__B2 (.I(\minimax.regD_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__I1 (.I(\minimax.regD_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__I1 (.I(\minimax.regD_uc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I1 (.I(\minimax.regD_uc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__I1 (.I(\minimax.regD_uc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I1 (.I(\minimax.regD_uc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__I1 (.I(\minimax.regD_uc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__A1 (.I(\minimax.regD_uc[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__A1 (.I(\minimax.regD_uc[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__I1 (.I(\minimax.regD_uc[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__I1 (.I(\minimax.regD_uc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__I1 (.I(\minimax.regD_uc[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__I1 (.I(\minimax.regD_uc[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__I1 (.I(\minimax.regD_uc[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__I1 (.I(\minimax.regD_uc[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__I1 (.I(\minimax.regD_uc[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__I1 (.I(\minimax.regD_uc[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I1 (.I(\minimax.regD_uc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__I1 (.I(\minimax.regD_uc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__I1 (.I(\minimax.regD_uc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__I1 (.I(\minimax.regD_uc[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__I1 (.I(\minimax.regD_uc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__I1 (.I(\minimax.regD_uc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(\minimax.regD_uc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__I1 (.I(\minimax.regD_uc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__I1 (.I(\minimax.regD_uc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__I1 (.I(\minimax.regD_uc[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__I1 (.I(\minimax.regD_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__I1 (.I(\minimax.regD_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__I1 (.I(\minimax.regD_uc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(\minimax.regD_uc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__I1 (.I(\minimax.regD_uc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I1 (.I(\minimax.regD_uc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__I1 (.I(\minimax.regD_uc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(\minimax.regD_uc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(\minimax.regD_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__I1 (.I(\minimax.regD_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(\minimax.regD_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__I1 (.I(\minimax.regD_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(\minimax.regD_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__I1 (.I(\minimax.regD_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A3 (.I(\minimax.regS_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(\minimax.regS_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A2 (.I(\minimax.regS_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__C (.I(\minimax.regS_ex[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(\minimax.regS_ex[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A2 (.I(\minimax.regS_ex[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(\minimax.regS_ex[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(\minimax.regS_ex[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I0 (.I(\minimax.regS_ex[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__I (.I(\minimax.regS_ex[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(\minimax.regS_ex[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(\minimax.regS_ex[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__I (.I(\minimax.regS_ex[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(\minimax.regS_ex[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A2 (.I(\minimax.regS_ex[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__I0 (.I(\minimax.regS_ex[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(\minimax.regS_ex[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A1 (.I(\minimax.regS_ex[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A3 (.I(\minimax.regS_ex[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__A1 (.I(\minimax.regS_ex[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A4 (.I(\minimax.regS_ex[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(\minimax.regS_ex[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(\minimax.regS_ex[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(\minimax.regS_ex[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(\minimax.regS_ex[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__I (.I(\minimax.regS_ex[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(\minimax.regS_ex[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(\minimax.regS_ex[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(\minimax.regS_ex[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(\minimax.regS_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__I (.I(\minimax.regS_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__C (.I(\minimax.regS_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(\minimax.regS_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B (.I(\minimax.regS_ex[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(\minimax.regS_ex[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(\minimax.regS_ex[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A3 (.I(\minimax.regS_ex[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__I (.I(\minimax.regS_ex[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__A1 (.I(\minimax.regS_ex[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(\minimax.regS_ex[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(\minimax.regS_ex[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A4 (.I(\minimax.regS_ex[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A1 (.I(\minimax.regS_ex[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(\minimax.regS_ex[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(\minimax.regS_ex[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(\minimax.regS_ex[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A3 (.I(\minimax.regS_ex[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A1 (.I(\minimax.regS_ex[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A2 (.I(\minimax.regS_ex[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(\minimax.regS_ex[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A4 (.I(\minimax.regS_ex[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A2 (.I(\minimax.regS_ex[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(\minimax.regS_ex[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(\minimax.regS_ex[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(\minimax.regS_ex[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A3 (.I(\minimax.regS_ex[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I0 (.I(\minimax.regS_ex[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A4 (.I(\minimax.regS_ex[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(\minimax.regS_ex[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(\minimax.regS_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(\minimax.regS_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__C (.I(\minimax.regS_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__B (.I(\minimax.regS_ex[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(\minimax.regS_ex[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I0 (.I(\minimax.regS_ex[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A3 (.I(\minimax.regS_ex[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(\minimax.regS_ex[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(\minimax.regS_ex[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__I (.I(\minimax.regS_ex[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__C (.I(\minimax.regS_ex[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I0 (.I(\minimax.regS_ex[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(\minimax.regS_ex[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(\minimax.regS_ex[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(\minimax.regS_ex[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(\minimax.regS_ex[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(\minimax.regS_ex[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(\minimax.regS_ex[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__B (.I(\minimax.regS_ex[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A3 (.I(\minimax.regS_ex[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__B (.I(\minimax.regS_ex[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__I (.I(\minimax.regS_ex[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A4 (.I(\minimax.regS_ex[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__I (.I(\minimax.regS_ex[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(\minimax.regS_ex[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(\minimax.regS_ex[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A3 (.I(\minimax.regS_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(\minimax.regS_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(\minimax.regS_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(\minimax.regS_uc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(\minimax.regS_uc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A2 (.I(\minimax.regS_uc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A1 (.I(\minimax.regS_uc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A1 (.I(\minimax.regS_uc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__I1 (.I(\minimax.regS_uc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__I (.I(\minimax.regS_uc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(\minimax.regS_uc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(\minimax.regS_uc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__A1 (.I(\minimax.regS_uc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__I (.I(\minimax.regS_uc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A2 (.I(\minimax.regS_uc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(\minimax.regS_uc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__I1 (.I(\minimax.regS_uc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(\minimax.regS_uc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(\minimax.regS_uc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(\minimax.regS_uc[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(\minimax.regS_uc[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A3 (.I(\minimax.regS_uc[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(\minimax.regS_uc[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(\minimax.regS_uc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(\minimax.regS_uc[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A3 (.I(\minimax.regS_uc[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__I (.I(\minimax.regS_uc[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(\minimax.regS_uc[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A1 (.I(\minimax.regS_uc[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A1 (.I(\minimax.regS_uc[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(\minimax.regS_uc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(\minimax.regS_uc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__I0 (.I(\minimax.regS_uc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__B (.I(\minimax.regS_uc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(\minimax.regS_uc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A2 (.I(\minimax.regS_uc[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A1 (.I(\minimax.regS_uc[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A4 (.I(\minimax.regS_uc[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__I (.I(\minimax.regS_uc[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(\minimax.regS_uc[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\minimax.regS_uc[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A1 (.I(\minimax.regS_uc[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A4 (.I(\minimax.regS_uc[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(\minimax.regS_uc[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(\minimax.regS_uc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A1 (.I(\minimax.regS_uc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A1 (.I(\minimax.regS_uc[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A3 (.I(\minimax.regS_uc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(\minimax.regS_uc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(\minimax.regS_uc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(\minimax.regS_uc[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A4 (.I(\minimax.regS_uc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(\minimax.regS_uc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(\minimax.regS_uc[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(\minimax.regS_uc[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A1 (.I(\minimax.regS_uc[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A3 (.I(\minimax.regS_uc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I1 (.I(\minimax.regS_uc[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A4 (.I(\minimax.regS_uc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(\minimax.regS_uc[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(\minimax.regS_uc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__I (.I(\minimax.regS_uc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(\minimax.regS_uc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I1 (.I(\minimax.regS_uc[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A3 (.I(\minimax.regS_uc[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(\minimax.regS_uc[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(\minimax.regS_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__I (.I(\minimax.regS_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__C (.I(\minimax.regS_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B (.I(\minimax.regS_uc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I1 (.I(\minimax.regS_uc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(\minimax.regS_uc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(\minimax.regS_uc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A1 (.I(\minimax.regS_uc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(\minimax.regS_uc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A1 (.I(\minimax.regS_uc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(\minimax.regS_uc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__B (.I(\minimax.regS_uc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A1 (.I(\minimax.regS_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A3 (.I(\minimax.regS_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(\minimax.regS_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__B (.I(\minimax.regS_uc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A1 (.I(\minimax.regS_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A4 (.I(\minimax.regS_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(\minimax.regS_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(\minimax.regS_uc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A1 (.I(\minimax.regS_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(\minimax.regS_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__A1 (.I(\minimax.regS_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(\minimax.regS_uc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2851__A3 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3565__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__A2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__I0 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__I0 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__I0 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__I0 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__I0 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__I0 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__I0 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__I1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__I1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__I1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__I1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__I0 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__I1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output86_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__I1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output87_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A2 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output88_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__I1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output89_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__I1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__I1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__I1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__I1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__I0 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__I1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__I1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__I0 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I0 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I0 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__I0 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__I0 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__I0 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[6]  (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[6]  (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[6]  (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[6]  (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[6]  (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[6]  (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[6]  (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[6]  (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[6]  (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[6]  (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[6]  (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[6]  (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[6]  (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[6]  (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[6]  (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[6]  (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[5]  (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[5]  (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[5]  (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[5]  (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[5]  (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[5]  (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[5]  (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[5]  (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[5]  (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[5]  (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[5]  (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[5]  (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[5]  (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[5]  (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[5]  (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[5]  (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[3]  (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[3]  (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[3]  (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[3]  (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[3]  (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[3]  (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[3]  (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[3]  (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[3]  (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[3]  (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[3]  (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[3]  (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[3]  (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[3]  (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[3]  (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[3]  (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[8]  (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[8]  (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[8]  (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[8]  (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[8]  (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[8]  (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[8]  (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[8]  (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[8]  (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[8]  (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[8]  (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[8]  (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[8]  (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[8]  (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[8]  (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[8]  (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[7]  (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[7]  (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[7]  (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[7]  (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[7]  (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[7]  (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[7]  (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[7]  (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[7]  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[7]  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[7]  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[7]  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[7]  (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[7]  (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[7]  (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[7]  (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[2]  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[2]  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[2]  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[2]  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[2]  (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[2]  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[2]  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[2]  (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[2]  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[2]  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[2]  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[2]  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[2]  (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[2]  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[2]  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[2]  (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[4]  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[4]  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[4]  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[4]  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[4]  (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[4]  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[4]  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[4]  (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[4]  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[4]  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[4]  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[4]  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[4]  (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[4]  (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[4]  (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[4]  (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[1]  (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[1]  (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[1]  (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[1]  (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[1]  (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[1]  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[1]  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[1]  (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[1]  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[1]  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[1]  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[1]  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[1]  (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[1]  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[1]  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[1]  (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_A[0]  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_A[0]  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_A[0]  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_A[0]  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_A[0]  (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_A[0]  (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_A[0]  (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_A[0]  (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_A[0]  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_A[0]  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_A[0]  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_A[0]  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_A[0]  (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_A[0]  (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_A[0]  (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_A[0]  (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram4_GWEN  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram1_GWEN  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram2_GWEN  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram1_GWEN  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram2_GWEN  (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram3_GWEN  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank1.ram4_GWEN  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank2.ram3_GWEN  (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram1_GWEN  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram2_GWEN  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram1_GWEN  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram2_GWEN  (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram3_GWEN  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank3.ram4_GWEN  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram3_GWEN  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_bank4.ram4_GWEN  (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout166_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer24_I (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__B (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__B (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A3 (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A4 (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer32_I (.I(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__B2 (.I(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__A4 (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A3 (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__A3 (.I(net397));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer48_I (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__I (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A3 (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_259_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_263_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_267_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_267_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_269_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_269_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_271_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_271_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_273_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_273_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_275_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_275_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_277_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_277_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_279_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_279_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_281_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_281_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_282_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_282_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_283_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_283_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_285_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_285_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_287_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_287_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_289_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_289_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_291_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_291_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_293_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_293_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_295_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_295_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_296_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_296_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_297_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_297_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_299_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_299_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_301_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_301_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_302_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_302_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_303_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_303_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_305_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_305_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_307_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_307_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_308_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_308_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_309_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_309_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_311_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_311_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_313_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_313_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_315_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_315_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_317_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_317_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_318_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_318_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_319_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_319_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_321_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_321_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_323_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_323_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_325_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_325_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_327_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_327_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_328_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_328_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_328_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_329_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_329_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_329_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_329_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_330_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_330_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_330_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_330_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_331_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_331_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_331_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_331_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_331_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_331_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_331_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_331_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_331_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_332_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_332_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_332_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_333_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_333_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_333_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_333_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_334_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_334_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_335_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_335_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_335_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_335_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_336_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_336_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_336_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_336_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_338_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_338_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_338_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_338_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_339_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_339_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_339_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_339_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_340_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_340_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_340_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_340_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_341_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_341_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_341_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_341_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_342_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_342_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_342_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_342_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_343_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_343_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_343_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_343_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_344_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_344_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_344_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_344_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_346_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_346_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_346_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_346_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_347_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_347_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_347_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_347_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_348_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_348_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_349_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_349_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_349_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_349_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_351_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_351_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_351_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_351_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_351_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_351_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_351_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_351_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_352_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_352_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_352_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_352_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_353_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_353_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_353_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_353_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_353_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_353_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_353_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_353_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_354_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_354_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_354_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_354_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_355_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_355_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_355_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_355_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_355_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_355_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_355_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_355_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_356_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_356_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_356_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_356_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_357_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_357_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_357_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_357_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_357_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_357_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_357_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_357_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_358_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_358_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_358_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_358_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_359_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_359_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_359_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_359_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_359_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_359_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_359_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_359_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_360_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_360_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_360_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_360_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_361_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_361_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_361_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_361_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_361_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_361_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_361_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_361_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_362_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_362_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_362_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_362_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_363_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_363_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_363_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_363_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_363_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_363_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_363_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_363_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_364_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_364_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_364_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_364_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_365_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_365_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_365_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_365_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_365_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_365_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_365_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_365_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_366_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_366_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_366_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_366_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_367_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_367_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_367_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_367_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_367_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_367_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_367_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_367_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_368_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_368_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_368_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_368_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_369_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_369_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_369_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_369_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_369_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_369_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_369_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_369_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_370_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_370_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_370_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_370_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_371_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_371_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_371_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_371_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_371_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_372_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_373_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_374_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_374_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_374_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_374_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_374_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_375_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_375_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_375_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_375_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_375_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_375_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_375_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_376_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_376_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_376_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_376_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_376_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_377_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_377_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_377_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_377_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_377_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_377_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_377_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_378_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_378_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_378_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_378_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_378_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_378_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_378_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_378_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_378_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_378_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_378_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_378_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_379_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_379_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_379_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_379_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_379_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_379_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_379_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_379_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_379_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_379_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_379_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_379_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_379_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_379_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_379_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_380_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_380_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_380_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_380_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_380_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_380_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_380_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_380_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_380_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_380_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_381_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_381_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_381_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_381_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_381_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_381_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_381_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_381_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_381_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_381_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_381_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_381_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_381_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_381_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_381_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_382_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_382_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_382_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_382_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_382_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_382_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_382_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_382_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_382_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_382_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_382_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_382_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_383_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_383_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_383_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_383_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_383_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_383_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_383_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_383_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_383_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_383_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_383_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_383_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_383_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_383_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_383_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_384_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_384_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_384_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_384_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_384_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_384_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_384_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_384_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_384_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_384_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_384_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_384_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_385_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_385_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_385_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_385_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_385_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_385_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_385_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_385_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_385_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_385_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_385_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_385_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_385_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_385_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_385_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_386_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_386_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_386_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_386_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_386_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_386_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_386_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_386_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_386_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_386_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_386_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_386_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_387_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_387_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_387_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_387_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_387_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_387_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_387_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_387_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_387_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_387_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_387_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_387_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_387_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_387_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_387_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_388_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_388_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_388_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_388_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_388_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_388_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_388_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_388_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_388_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_388_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_388_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_388_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_389_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_389_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_389_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_389_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_389_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_389_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_389_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_389_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_389_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_389_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_389_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_389_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_389_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_389_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_389_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_390_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_390_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_390_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_390_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_390_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_390_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_390_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_390_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_390_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_390_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_391_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_391_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_391_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_391_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_391_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_391_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_391_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_391_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_391_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_391_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_391_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_391_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_391_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_391_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_391_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_392_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_392_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_392_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_392_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_392_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_392_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_392_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_392_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_392_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_392_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_392_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_392_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_393_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_393_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_393_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_393_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_393_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_393_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_393_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_393_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_393_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_393_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_393_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_393_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_393_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_393_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_393_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_394_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_394_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_394_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_394_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_394_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_394_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_394_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_394_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_394_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_394_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_394_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_394_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_395_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_395_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_395_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_395_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_395_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_395_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_395_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_395_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_395_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_395_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_395_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_395_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_395_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_395_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_395_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_396_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_396_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_396_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_396_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_396_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_396_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_396_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_396_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_396_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_396_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_396_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_396_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_397_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_397_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_397_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_397_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_397_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_397_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_397_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_397_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_397_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_397_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_397_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_397_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_397_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_397_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_397_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_398_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_398_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_398_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_398_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_398_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_398_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_398_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_398_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_398_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_398_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_398_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_398_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_399_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_399_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_399_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_399_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_399_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_399_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_399_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_399_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_399_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_399_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_399_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_399_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_399_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_399_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_399_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_400_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_400_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_400_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_400_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_400_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_400_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_400_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_400_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_400_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_400_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_401_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_401_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_401_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_401_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_401_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_401_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_401_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_401_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_401_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_401_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_401_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_401_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_401_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_401_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_401_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_402_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_402_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_402_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_402_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_402_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_402_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_402_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_402_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_402_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_402_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_402_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_402_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_403_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_403_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_403_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_403_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_403_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_403_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_403_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_403_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_403_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_403_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_403_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_403_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_403_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_403_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_403_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_404_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_404_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_404_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_404_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_404_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_404_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_404_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_404_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_404_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_404_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_404_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_404_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_405_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_405_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_405_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_405_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_405_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_405_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_405_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_405_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_405_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_405_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_405_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_405_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_405_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_405_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_405_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_406_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_406_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_406_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_406_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_406_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_406_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_406_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_406_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_406_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_406_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_406_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_406_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_407_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_407_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_407_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_407_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_407_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_407_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_407_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_407_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_407_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_407_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_407_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_407_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_407_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_407_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_407_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_408_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_408_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_408_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_408_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_408_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_408_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_408_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_408_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_408_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_408_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_408_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_408_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_409_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_409_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_409_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_409_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_409_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_409_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_409_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_409_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_409_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_409_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_409_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_409_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_409_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_409_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_409_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_410_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_410_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_410_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_410_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_410_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_410_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_410_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_410_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_410_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_410_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_410_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_410_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_411_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_411_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_411_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_411_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_411_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_411_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_411_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_411_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_411_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_411_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_411_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_411_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_411_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_412_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_412_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_412_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_412_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_412_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_412_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_412_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_412_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_412_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_412_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_412_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_412_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_413_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_413_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_413_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_413_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_413_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_413_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_413_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_413_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_413_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_413_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_413_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_413_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_413_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_413_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_413_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_414_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_414_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_414_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_414_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_414_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_414_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_414_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_414_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_414_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_414_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_414_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_414_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_415_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_415_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_415_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_415_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_415_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_415_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_415_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_415_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_415_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_415_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_415_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_415_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_415_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_415_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_415_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_416_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_416_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_416_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_416_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_416_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_416_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_416_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_416_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_416_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_416_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_416_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_416_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_417_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_417_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_417_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_417_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_417_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_417_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_417_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_417_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_417_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_417_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_417_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_417_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_417_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_417_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_417_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_418_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_418_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_418_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_418_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_418_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_418_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_418_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_418_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_418_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_418_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_418_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_418_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_419_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_419_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_419_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_419_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_419_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_419_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_419_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_419_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_419_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_419_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_419_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_419_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_419_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_419_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_420_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_420_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_420_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_420_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_420_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_420_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_420_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_420_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_420_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_421_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_421_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_421_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_421_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_421_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_421_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_421_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_421_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_421_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_421_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_422_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_422_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_422_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_422_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_422_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_422_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_422_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_422_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_422_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_423_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_423_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_423_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_423_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_423_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_423_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_423_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_424_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_424_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_424_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_424_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_424_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_424_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_424_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_425_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_425_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_425_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_425_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_425_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_425_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_425_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_425_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_425_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_425_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_425_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_425_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_425_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_425_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_425_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_426_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_426_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_426_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_426_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_426_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_426_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_426_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_426_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_426_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_426_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_426_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_426_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_427_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_427_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_427_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_427_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_427_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_427_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_427_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_427_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_427_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_427_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_427_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_427_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_427_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_427_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_427_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_427_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_427_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_427_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_428_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_428_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_428_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_428_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_428_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_428_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_428_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_428_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_428_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_428_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_428_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_428_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_429_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_429_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_429_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_429_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_429_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_429_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_429_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_429_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_429_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_429_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_429_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_429_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_429_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_429_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_429_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_430_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_430_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_430_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_430_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_430_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_430_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_430_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_430_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_430_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_430_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_430_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_430_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_431_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_431_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_431_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_431_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_431_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_431_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_431_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_431_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_431_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_431_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_431_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_431_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_431_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_431_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_431_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_431_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_431_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_432_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_432_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_432_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_432_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_432_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_432_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_432_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_432_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_432_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_432_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_432_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_432_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_433_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_433_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_433_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_433_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_433_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_433_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_433_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_433_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_433_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_433_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_433_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_433_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_433_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_433_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_433_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_434_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_434_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_434_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_434_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_434_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_434_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_434_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_434_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_434_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_434_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_434_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_434_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_435_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_435_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_435_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_435_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_435_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_435_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_435_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_435_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_435_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_435_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_435_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_435_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_435_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_435_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_435_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_436_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_436_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_436_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_436_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_436_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_436_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_436_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_436_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_436_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_436_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_436_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_436_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_437_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_437_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_437_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_437_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_437_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_437_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_437_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_437_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_437_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_437_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_437_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_437_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_437_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_437_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_437_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_438_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_438_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_438_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_438_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_438_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_438_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_438_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_438_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_438_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_438_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_438_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_438_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_439_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_439_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_439_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_439_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_439_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_439_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_439_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_439_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_439_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_439_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_439_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_439_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_439_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_439_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_439_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_439_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_439_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_439_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_440_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_440_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_440_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_440_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_440_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_440_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_440_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_440_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_440_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_440_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_440_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_440_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_441_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_441_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_441_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_441_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_441_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_441_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_441_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_441_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_441_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_441_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_441_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_441_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_441_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_441_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_441_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_441_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_441_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_442_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_442_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_442_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_442_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_442_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_442_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_442_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_442_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_442_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_442_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_442_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_442_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_443_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_443_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_443_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_443_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_443_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_443_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_443_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_443_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_443_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_443_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_443_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_443_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_443_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_443_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_443_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_444_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_444_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_444_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_444_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_444_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_444_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_444_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_444_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_444_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_444_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_444_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_444_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_445_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_445_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_445_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_445_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_445_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_445_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_445_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_445_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_445_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_445_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_445_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_445_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_445_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_445_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_445_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_446_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_446_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_446_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_446_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_446_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_446_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_446_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_446_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_446_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_446_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_446_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_446_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_447_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_447_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_447_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_447_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_447_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_447_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_447_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_447_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_447_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_447_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_447_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_447_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_447_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_447_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_447_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_447_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_447_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_447_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_448_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_448_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_448_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_448_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_448_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_448_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_448_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_448_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_448_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_448_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_448_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_448_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_449_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_449_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_449_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_449_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_449_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_449_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_449_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_449_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_449_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_449_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_449_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_449_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_449_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_449_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_449_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_449_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_449_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_449_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_450_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_450_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_450_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_450_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_450_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_450_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_450_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_450_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_450_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_450_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_450_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_450_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_451_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_451_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_451_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_451_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_451_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_451_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_451_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_451_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_451_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_451_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_451_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_451_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_451_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_451_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_451_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_451_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_451_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_451_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_451_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_451_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_452_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_452_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_452_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_452_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_452_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_452_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_452_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_452_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_452_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_452_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_452_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_452_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_453_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_453_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_453_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_453_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_453_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_453_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_453_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_453_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_453_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_453_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_453_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_453_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_453_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_453_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_453_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_453_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_453_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_453_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_454_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_454_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_454_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_454_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_454_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_454_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_454_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_454_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_454_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_454_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_454_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_454_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_455_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_455_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_455_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_455_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_455_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_455_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_455_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_455_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_455_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_455_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_455_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_455_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_455_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_455_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_455_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_456_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_456_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_456_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_456_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_456_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_456_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_456_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_456_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_456_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_456_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_456_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_456_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_457_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_457_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_457_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_457_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_457_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_457_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_457_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_457_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_457_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_457_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_457_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_457_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_457_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_457_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_457_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_458_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_458_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_458_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_458_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_458_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_458_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_458_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_458_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_458_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_458_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_458_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_458_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_459_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_459_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_459_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_459_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_459_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_459_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_459_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_459_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_459_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_459_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_459_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_459_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_459_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_459_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_459_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_460_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_460_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_460_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_460_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_460_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_460_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_460_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_460_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_460_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_460_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_460_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_460_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_461_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_461_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_461_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_461_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_461_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_461_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_461_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_461_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_461_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_461_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_461_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_461_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_461_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_461_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_461_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_461_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_461_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_462_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_462_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_462_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_462_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_462_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_462_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_462_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_462_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_462_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_462_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_462_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_462_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_463_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_463_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_463_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_463_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_463_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_463_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_463_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_463_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_463_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_463_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_463_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_463_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_463_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_463_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_463_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_464_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_464_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_464_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_464_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_464_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_464_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_464_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_464_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_464_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_464_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_464_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_464_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_465_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_465_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_465_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_465_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_465_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_465_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_465_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_465_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_465_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_465_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_465_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_465_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_465_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_465_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_465_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_466_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_466_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_466_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_466_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_466_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_466_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_466_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_466_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_466_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_466_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_466_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_466_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_467_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_467_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_467_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_467_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_467_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_467_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_467_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_467_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_467_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_467_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_467_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_467_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_467_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_467_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_467_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_468_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_468_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_468_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_468_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_468_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_468_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_468_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_468_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_468_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_468_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_468_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_468_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_469_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_469_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_469_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_469_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_469_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_469_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_469_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_469_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_469_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_469_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_469_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_469_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_469_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_469_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_469_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_470_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_470_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_470_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_470_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_470_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_470_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_470_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_470_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_470_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_470_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_470_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_470_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_471_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_471_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_471_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_471_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_471_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_471_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_471_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_471_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_471_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_471_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_471_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_471_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_471_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_471_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_471_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_471_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_471_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_472_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_472_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_472_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_472_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_472_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_472_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_472_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_472_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_472_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_472_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_472_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_472_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_473_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_473_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_473_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_473_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_473_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_473_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_473_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_473_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_473_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_473_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_473_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_473_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_473_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_473_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_473_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_474_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_474_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_474_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_474_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_474_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_474_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_474_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_474_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_474_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_474_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_474_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_474_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_475_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_475_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_475_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_475_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_475_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_475_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_475_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_475_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_475_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_475_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_475_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_475_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_475_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_475_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_475_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_476_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_476_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_476_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_476_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_476_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_476_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_476_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_476_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_476_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_476_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_476_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_476_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_477_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_477_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_477_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_477_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_477_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_477_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_477_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_477_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_477_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_477_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_477_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_477_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_477_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_477_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_477_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_478_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_478_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_478_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_478_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_478_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_478_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_478_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_478_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_478_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_478_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_478_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_478_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_479_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_479_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_479_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_479_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_479_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_479_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_479_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_479_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_479_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_479_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_479_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_479_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_479_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_479_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_479_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_480_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_480_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_480_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_480_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_480_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_480_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_480_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_480_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_480_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_480_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_480_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_480_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_481_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_481_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_481_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_481_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_481_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_481_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_481_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_481_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_481_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_481_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_481_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_481_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_481_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_481_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_481_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_482_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_482_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_482_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_482_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_482_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_482_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_482_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_482_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_482_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_482_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_482_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_482_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_482_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_482_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_482_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_482_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_482_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_483_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_483_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_483_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_483_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_483_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_483_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_483_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_483_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_483_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_483_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_483_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_483_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_483_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_483_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_483_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_484_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_484_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_484_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_484_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_484_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_484_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_484_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_484_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_484_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_484_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_484_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_484_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_485_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_485_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_485_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_485_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_485_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_485_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_485_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_485_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_485_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_485_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_485_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_485_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_485_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_485_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_485_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_486_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_486_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_486_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_486_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_486_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_486_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_486_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_486_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_486_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_486_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_486_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_486_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_487_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_487_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_487_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_487_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_487_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_487_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_487_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_487_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_487_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_487_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_487_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_487_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_487_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_487_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_487_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_488_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_488_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_488_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_488_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_488_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_488_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_488_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_488_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_488_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_488_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_488_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_488_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_489_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_489_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_489_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_489_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_489_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_489_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_489_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_489_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_489_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_489_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_489_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_489_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_489_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_489_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_489_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_490_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_490_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_490_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_490_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_490_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_490_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_491_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_491_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_491_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_491_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_491_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_491_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_491_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_491_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_491_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_491_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_491_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_491_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_491_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_491_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_492_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_492_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_492_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_492_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_492_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_492_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_492_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_492_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_492_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_492_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_493_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_493_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_493_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_493_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_493_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_493_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_493_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_493_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_493_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_493_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_493_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_493_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_493_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_493_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_494_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_494_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_494_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_495_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_495_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_495_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_496_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_496_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_496_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_496_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_496_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_496_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_497_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_497_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_497_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_498_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_498_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_498_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_498_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_498_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_498_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_499_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_499_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_499_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_499_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_499_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_499_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_499_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_499_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_499_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_499_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_499_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_499_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_499_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_500_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_500_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_500_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_500_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_500_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_500_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_500_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_501_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_501_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_501_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_501_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_501_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_501_5330 ();
 assign io_oeb[37] = net169;
 assign io_out[0] = net170;
 assign io_out[10] = net180;
 assign io_out[11] = net181;
 assign io_out[12] = net182;
 assign io_out[13] = net183;
 assign io_out[14] = net184;
 assign io_out[15] = net185;
 assign io_out[16] = net186;
 assign io_out[17] = net187;
 assign io_out[18] = net188;
 assign io_out[19] = net189;
 assign io_out[1] = net171;
 assign io_out[20] = net190;
 assign io_out[21] = net191;
 assign io_out[22] = net192;
 assign io_out[23] = net193;
 assign io_out[24] = net194;
 assign io_out[25] = net195;
 assign io_out[26] = net196;
 assign io_out[27] = net197;
 assign io_out[28] = net198;
 assign io_out[29] = net199;
 assign io_out[2] = net172;
 assign io_out[30] = net200;
 assign io_out[31] = net201;
 assign io_out[32] = net202;
 assign io_out[33] = net203;
 assign io_out[34] = net204;
 assign io_out[35] = net205;
 assign io_out[36] = net206;
 assign io_out[37] = net207;
 assign io_out[3] = net173;
 assign io_out[4] = net174;
 assign io_out[5] = net175;
 assign io_out[6] = net176;
 assign io_out[7] = net177;
 assign io_out[8] = net178;
 assign io_out[9] = net179;
 assign irq[0] = net208;
 assign irq[1] = net209;
 assign irq[2] = net210;
 assign la_data_out[0] = net211;
 assign la_data_out[100] = net311;
 assign la_data_out[101] = net312;
 assign la_data_out[102] = net313;
 assign la_data_out[103] = net314;
 assign la_data_out[104] = net315;
 assign la_data_out[105] = net316;
 assign la_data_out[106] = net317;
 assign la_data_out[107] = net318;
 assign la_data_out[108] = net319;
 assign la_data_out[109] = net320;
 assign la_data_out[10] = net221;
 assign la_data_out[110] = net321;
 assign la_data_out[111] = net322;
 assign la_data_out[112] = net323;
 assign la_data_out[113] = net324;
 assign la_data_out[114] = net325;
 assign la_data_out[115] = net326;
 assign la_data_out[116] = net327;
 assign la_data_out[117] = net328;
 assign la_data_out[118] = net329;
 assign la_data_out[119] = net330;
 assign la_data_out[11] = net222;
 assign la_data_out[120] = net331;
 assign la_data_out[121] = net332;
 assign la_data_out[122] = net333;
 assign la_data_out[123] = net334;
 assign la_data_out[124] = net335;
 assign la_data_out[125] = net336;
 assign la_data_out[126] = net337;
 assign la_data_out[127] = net338;
 assign la_data_out[12] = net223;
 assign la_data_out[13] = net224;
 assign la_data_out[14] = net225;
 assign la_data_out[15] = net226;
 assign la_data_out[16] = net227;
 assign la_data_out[17] = net228;
 assign la_data_out[18] = net229;
 assign la_data_out[19] = net230;
 assign la_data_out[1] = net212;
 assign la_data_out[20] = net231;
 assign la_data_out[21] = net232;
 assign la_data_out[22] = net233;
 assign la_data_out[23] = net234;
 assign la_data_out[24] = net235;
 assign la_data_out[25] = net236;
 assign la_data_out[26] = net237;
 assign la_data_out[27] = net238;
 assign la_data_out[28] = net239;
 assign la_data_out[29] = net240;
 assign la_data_out[2] = net213;
 assign la_data_out[30] = net241;
 assign la_data_out[31] = net242;
 assign la_data_out[32] = net243;
 assign la_data_out[33] = net244;
 assign la_data_out[34] = net245;
 assign la_data_out[35] = net246;
 assign la_data_out[36] = net247;
 assign la_data_out[37] = net248;
 assign la_data_out[38] = net249;
 assign la_data_out[39] = net250;
 assign la_data_out[3] = net214;
 assign la_data_out[40] = net251;
 assign la_data_out[41] = net252;
 assign la_data_out[42] = net253;
 assign la_data_out[43] = net254;
 assign la_data_out[44] = net255;
 assign la_data_out[45] = net256;
 assign la_data_out[46] = net257;
 assign la_data_out[47] = net258;
 assign la_data_out[48] = net259;
 assign la_data_out[49] = net260;
 assign la_data_out[4] = net215;
 assign la_data_out[50] = net261;
 assign la_data_out[51] = net262;
 assign la_data_out[52] = net263;
 assign la_data_out[53] = net264;
 assign la_data_out[54] = net265;
 assign la_data_out[55] = net266;
 assign la_data_out[56] = net267;
 assign la_data_out[57] = net268;
 assign la_data_out[58] = net269;
 assign la_data_out[59] = net270;
 assign la_data_out[5] = net216;
 assign la_data_out[60] = net271;
 assign la_data_out[61] = net272;
 assign la_data_out[62] = net273;
 assign la_data_out[63] = net274;
 assign la_data_out[64] = net275;
 assign la_data_out[65] = net276;
 assign la_data_out[66] = net277;
 assign la_data_out[67] = net278;
 assign la_data_out[68] = net279;
 assign la_data_out[69] = net280;
 assign la_data_out[6] = net217;
 assign la_data_out[70] = net281;
 assign la_data_out[71] = net282;
 assign la_data_out[72] = net283;
 assign la_data_out[73] = net284;
 assign la_data_out[74] = net285;
 assign la_data_out[75] = net286;
 assign la_data_out[76] = net287;
 assign la_data_out[77] = net288;
 assign la_data_out[78] = net289;
 assign la_data_out[79] = net290;
 assign la_data_out[7] = net218;
 assign la_data_out[80] = net291;
 assign la_data_out[81] = net292;
 assign la_data_out[82] = net293;
 assign la_data_out[83] = net294;
 assign la_data_out[84] = net295;
 assign la_data_out[85] = net296;
 assign la_data_out[86] = net297;
 assign la_data_out[87] = net298;
 assign la_data_out[88] = net299;
 assign la_data_out[89] = net300;
 assign la_data_out[8] = net219;
 assign la_data_out[90] = net301;
 assign la_data_out[91] = net302;
 assign la_data_out[92] = net303;
 assign la_data_out[93] = net304;
 assign la_data_out[94] = net305;
 assign la_data_out[95] = net306;
 assign la_data_out[96] = net307;
 assign la_data_out[97] = net308;
 assign la_data_out[98] = net309;
 assign la_data_out[99] = net310;
 assign la_data_out[9] = net220;
 assign wbs_ack_o = net339;
endmodule

