module minimax (clk,
    inst_regce,
    reset,
    rreq,
    vdd,
    vss,
    wb,
    addr,
    addrD,
    addrS,
    aluX,
    inst,
    inst_addr,
    rdata,
    regD,
    regS,
    wdata,
    wmask);
 input clk;
 output inst_regce;
 input reset;
 output rreq;
 input vdd;
 input vss;
 output wb;
 output [31:0] addr;
 output [5:0] addrD;
 output [5:0] addrS;
 output [31:0] aluX;
 input [15:0] inst;
 output [11:0] inst_addr;
 input [31:0] rdata;
 input [31:0] regD;
 input [31:0] regS;
 output [31:0] wdata;
 output [3:0] wmask;

 wire net147;
 wire net173;
 wire net162;
 wire net161;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net155;
 wire net154;
 wire net153;
 wire net152;
 wire net172;
 wire net151;
 wire net150;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire net171;
 wire net160;
 wire net170;
 wire net149;
 wire net148;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire bubble1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A3;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A2;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN;
 wire bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1;
 wire bubble2;
 wire bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire dly16_lw;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN;
 wire dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN;
 wire dly16_lwsp;
 wire dly16_slli_setrd;
 wire dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1;
 wire dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3;
 wire dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN;
 wire dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2;
 wire dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z;
 wire dly16_slli_setrs;
 wire dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1;
 wire dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_A1;
 wire dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z;
 wire \dra[0] ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_ZN ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ;
 wire \dra[1] ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ;
 wire \dra[2] ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1 ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ;
 wire \dra[3] ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A4 ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ;
 wire \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ;
 wire \dra[4] ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ;
 wire \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ;
 wire inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D;
 wire microcode;
 wire microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN;
 wire microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D;
 wire microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2;
 wire microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire op16_lw;
 wire op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I;
 wire op16_lwsp;
 wire op16_slli_setrd;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_C;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_A2;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN;
 wire op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2;
 wire op16_slli_setrs;
 wire op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2;
 wire op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2;
 wire op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2;
 wire op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN;
 wire \pc_execute[10] ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ;
 wire \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[11] ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ;
 wire \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ;
 wire \pc_execute[1] ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ;
 wire \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ;
 wire \pc_execute[2] ;
 wire \pc_execute[3] ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A4 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ;
 wire \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_ZN ;
 wire \pc_execute[4] ;
 wire \pc_execute[5] ;
 wire \pc_execute[6] ;
 wire \pc_execute[7] ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ;
 wire \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ;
 wire \pc_execute[8] ;
 wire \pc_execute[9] ;
 wire \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_B ;
 wire \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ;
 wire \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ;
 wire \pc_fetch_dly[10] ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_fetch_dly[11] ;
 wire \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[1] ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ;
 wire \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_fetch_dly[2] ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ;
 wire \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire \pc_fetch_dly[3] ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_Z ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ;
 wire \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_fetch_dly[4] ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ;
 wire \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_fetch_dly[5] ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ;
 wire \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire \pc_fetch_dly[6] ;
 wire \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ;
 wire \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ;
 wire \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire \pc_fetch_dly[7] ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ;
 wire \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[8] ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ;
 wire \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ;
 wire \pc_fetch_dly[9] ;
 wire \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ;
 wire \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ;
 wire \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ;
 wire \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ;
 wire \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ;
 wire reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z;
 wire reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z;
 wire reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_A2;
 wire reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_ZN;
 wire wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I;
 wire wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_1_I (.I(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_3_I (.I(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_8_I (.I(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_9_I (.I(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A2 (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3 (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A3 (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_A3 (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_S (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 (.I(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 (.I(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__or2_2_A2_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__or2_2_A2_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z_I (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_B (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_4_Z_I (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A3 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D (.I(bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D (.I(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A1 (.I(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A1 (.I(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A1 (.I(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A1 (.I(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A1 (.I(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A1 (.I(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lwsp_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_lwsp_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D (.I(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A2 (.I(dly16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A1 (.I(dly16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A2 (.I(dly16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1 (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_1_A2 (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_1_B (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_2_A2 (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_2_B (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_A2 (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_B (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_A2 (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_B (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A2 (.I(dly16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I (.I(dly16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A2 (.I(dly16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_B2  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B  (.I(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2  (.I(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2  (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A1  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1  (.I(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_1_C_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_1_C_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_Z_I  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_2_ZN_A1  (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_2_ZN_A2  (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_2_ZN_A3  (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_2_ZN_A4  (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_I  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A1  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A2  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1  (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A3_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3  (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__inv_2_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_B  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A1  (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1  (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1  (.I(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A1  (.I(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A2  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I  (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2  (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_2_B_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_2_B_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A1  (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A2  (.I(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1  (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2  (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3  (.I(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_B  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B  (.I(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_B1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_B2  (.I(\dra[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A3  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_1_I_I  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\dra[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A2  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C  (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z_I  (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(inst[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(inst[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(inst[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(inst[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(inst[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(inst[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(inst[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(rdata[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(rdata[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(rdata[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(inst[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(rdata[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(rdata[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(rdata[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(rdata[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(rdata[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(rdata[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(rdata[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(rdata[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(rdata[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(rdata[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(inst[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(rdata[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(rdata[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(rdata[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(rdata[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(rdata[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(rdata[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(rdata[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(rdata[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(rdata[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(rdata[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(inst[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(rdata[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(rdata[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(rdata[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(rdata[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(rdata[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(rdata[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(rdata[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(rdata[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(rdata[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(reset),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(inst[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(inst[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(inst[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(inst[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(inst[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(inst[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D (.I(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z_I (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2 (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_C (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_lwsp_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1 (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_lwsp_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A2 (.I(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_D (.I(op16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A2 (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_B1 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_B2 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_B1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A2 (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 (.I(net135),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I0 (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_S (.I(\pc_execute[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_A1 (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 (.I(\pc_execute[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B2 (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I (.I(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A1 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_D (.I(op16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output90_I (.I(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output91_I (.I(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2  (.I(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_B  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_B  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\pc_execute[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_A2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3  (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_C  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_B  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_S  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(\pc_fetch_dly[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A4_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A4_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A4_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A4_A4  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1  (.I(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A2  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A2  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_execute[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(\pc_fetch_dly[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\pc_execute[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A2  (.I(\pc_execute[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A2  (.I(\pc_execute[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A1  (.I(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_B  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2  (.I(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z_I  (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN_A1  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN_B  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN_A1  (.I(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3  (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_A4  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_C  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2  (.I(\pc_execute[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A1  (.I(\pc_execute[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_B  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C  (.I(\pc_execute[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\pc_execute[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\pc_execute[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A3  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A4  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A1  (.I(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A1  (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(\pc_fetch_dly[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z_I  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1  (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(net134),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_2_A1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_B  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_1_A1  (.I(\pc_execute[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_1_B  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_A1  (.I(\pc_execute[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_A2  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1  (.I(net136),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\pc_fetch_dly[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\pc_fetch_dly[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\pc_fetch_dly[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1  (.I(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_A1  (.I(\pc_fetch_dly[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\pc_fetch_dly[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A1  (.I(\pc_fetch_dly[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B2  (.I(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C2  (.I(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I0  (.I(\pc_execute[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I1  (.I(\pc_fetch_dly[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_S  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\pc_fetch_dly[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I  (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I_I  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A1  (.I(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2  (.I(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_A1  (.I(\pc_fetch_dly[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\pc_fetch_dly[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\pc_fetch_dly[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I_I  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN_I  (.I(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I1  (.I(\pc_fetch_dly[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_S  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\pc_fetch_dly[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A1  (.I(\pc_fetch_dly[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1  (.I(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A1  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B2  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I_I  (.I(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I0  (.I(\pc_execute[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I1  (.I(\pc_fetch_dly[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_S  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B2  (.I(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C1  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C2  (.I(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I0  (.I(\pc_execute[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_S  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A1  (.I(\pc_fetch_dly[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A1  (.I(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A1  (.I(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A1  (.I(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A1  (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1  (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_4_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_4_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B2  (.I(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C1  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C2  (.I(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net134),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_A1  (.I(\pc_fetch_dly[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_B1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_B2  (.I(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_C1  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_C2  (.I(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I_I  (.I(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net135),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A1  (.I(\pc_fetch_dly[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2  (.I(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A1  (.I(\pc_fetch_dly[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B2  (.I(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C1  (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_C2  (.I(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I_I  (.I(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I0  (.I(\pc_fetch_dly[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_I1  (.I(net136),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I0  (.I(\pc_execute[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_I1  (.I(\pc_fetch_dly[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_S  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_I (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_A1 (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D_CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rreq_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A1 (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A2 (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3 (.I(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A1 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_B (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_1_I (.I(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_2_I (.I(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I (.I(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_13 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(net146),
    .Z(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_1 (.I(net78),
    .Z(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_10 (.I(net145),
    .Z(net85),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_2 (.I(net144),
    .Z(net75),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_3 (.I(net146),
    .Z(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_4 (.I(net144),
    .Z(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_5 (.I(net144),
    .Z(net79),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_6 (.I(net144),
    .Z(net80),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_7 (.I(net144),
    .Z(net81),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_8 (.I(net146),
    .Z(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 addr_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_9 (.I(net146),
    .Z(net83),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .CLK(clknet_2_1__leaf_clk),
    .Q(bubble1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z (.A1(bubble2),
    .A2(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .A3(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2 (.A1(bubble2),
    .A2(bubble1),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2 (.A1(bubble2),
    .A2(bubble1),
    .A3(net1),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2 (.A1(bubble2),
    .A2(bubble1),
    .A3(net1),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3),
    .ZN(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z (.A1(net7),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A3),
    .A4(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z (.I0(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3 ),
    .I1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I1),
    .S(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A2(net4),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A4_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z_I1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3 (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A2),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN),
    .A4(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .A4(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(net10),
    .A2(net9),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A4_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(net8),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_4_Z (.I(net6),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN (.I(net5),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S (.I0(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .I1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .S(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__or2_2_A2 (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2 (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_4_Z (.I(net7),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .CLK(clknet_2_1__leaf_clk),
    .Q(bubble2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .ZN(bubble2_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(op16_lw),
    .CLK(clknet_2_3__leaf_clk),
    .Q(dly16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2 (.A1(dly16_lwsp),
    .A2(dly16_lw),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z),
    .Z(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(net34),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1 (.A1(net33),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2 (.A1(net32),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3 (.A1(net31),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4 (.A1(net30),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(net29),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1 (.A1(net27),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2 (.A1(net26),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3 (.A1(net25),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3 (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .Z(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(net23),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1 (.A1(net22),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2 (.A1(net21),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3 (.A1(net20),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4 (.A1(net17),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(net40),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1 (.A1(net38),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2 (.A1(net37),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3 (.A1(net36),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4 (.A1(net35),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 dly16_lwsp_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(op16_lwsp),
    .CLK(clknet_2_3__leaf_clk),
    .Q(dly16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2 (.A1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(dly16_slli_setrd),
    .A3(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .ZN(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN),
    .A2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1 (.A1(dly16_slli_setrd),
    .A2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .Z(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2 (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN),
    .A2(dly16_slli_setrd),
    .Z(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .A2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z),
    .ZN(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2 (.A1(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .A2(dly16_slli_setrs),
    .B(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B (.A1(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .B(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .ZN(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_1 (.A1(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .B(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .ZN(net86),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_B_2 (.A1(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .B(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .ZN(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B (.A1(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_A1),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .B(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .ZN(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .Z(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(dly16_slli_setrs),
    .Z(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2 (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN),
    .A2(dly16_slli_setrs),
    .Z(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .A2(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z),
    .ZN(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1  (.A1(\dra[0] ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .C(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .Z(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_ZN ),
    .ZN(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\dra[0] ),
    .A2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .Z(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .Z(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .A2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .ZN(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .B(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net14),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\dra[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(op16_lw),
    .B1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B2(net14),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .A2(\dra[1] ),
    .B(op16_lwsp),
    .C(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .A2(op16_lwsp),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .B2(net14),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .A3(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .ZN(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net15),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A3(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3 ),
    .ZN(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(op16_lwsp),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .B(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A2_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_1_C  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .B(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .C(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ),
    .ZN(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\dra[1] ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .A3(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .ZN(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_Z  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2 ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2 ),
    .B(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_2_ZN  (.A1(net2),
    .A2(net3),
    .A3(net16),
    .A4(net14),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net15),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\dra[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(op16_lw),
    .B1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .ZN(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\dra[2] ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .A2(\dra[2] ),
    .B1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .Z(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .A2(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .B(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN ),
    .ZN(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net16),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .B1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1 ),
    .B2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .C(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .ZN(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .B(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\dra[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .A2(op16_lw),
    .B1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B2(net16),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .A2(\dra[3] ),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN  (.A1(net6),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A2(net4),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1_ZN ),
    .ZN(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(net13),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .Z(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_2_A3  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN  (.A1(net6),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .A3(net7),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .A4(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net2),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .ZN(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .Z(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__inv_2_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .ZN(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z  (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2  (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2  (.A1(net133),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3  (.A1(net132),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .A4(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(net4),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN  (.A1(net6),
    .A2(net7),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai211_2_B  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_ZN ),
    .C(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B2(\dra[3] ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_4_A2_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN ),
    .A4(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A4 ),
    .ZN(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN  (.A1(net3),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .B(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .A2(net9),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .A4(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN  (.A1(net13),
    .A2(net12),
    .A3(net11),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .Z(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net8),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\dra[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B(op16_lw),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .B1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B2(\dra[4] ),
    .C1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1 ),
    .C2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net2),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .A3(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_A3  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A3(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net3),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_1_I  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_ZN ),
    .ZN(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\dra[4] ),
    .A2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net13),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN),
    .C(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A3(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3 ),
    .A4(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and4_1_Z_A4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\dra[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ),
    .A3(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net3),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN_I_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z  (.I(net1),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .Z(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ),
    .Z(op16_lwsp),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout144 (.I(net145),
    .Z(net144),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net146),
    .Z(net145),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout146 (.I(net86),
    .Z(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input1 (.I(inst[0]),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(inst[3]),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(inst[4]),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(inst[5]),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(inst[6]),
    .Z(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input14 (.I(inst[7]),
    .Z(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input15 (.I(inst[8]),
    .Z(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input16 (.I(inst[9]),
    .Z(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(rdata[0]),
    .Z(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(rdata[10]),
    .Z(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(rdata[11]),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(inst[10]),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(rdata[12]),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(rdata[13]),
    .Z(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input22 (.I(rdata[14]),
    .Z(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(rdata[15]),
    .Z(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input24 (.I(rdata[16]),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(rdata[17]),
    .Z(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(rdata[18]),
    .Z(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(rdata[19]),
    .Z(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(rdata[1]),
    .Z(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(rdata[20]),
    .Z(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(inst[11]),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(rdata[21]),
    .Z(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(rdata[22]),
    .Z(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(rdata[23]),
    .Z(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(rdata[24]),
    .Z(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(rdata[25]),
    .Z(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(rdata[26]),
    .Z(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(rdata[27]),
    .Z(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(rdata[28]),
    .Z(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(rdata[29]),
    .Z(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input39 (.I(rdata[2]),
    .Z(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(inst[12]),
    .Z(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input40 (.I(rdata[30]),
    .Z(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(rdata[31]),
    .Z(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(rdata[3]),
    .Z(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input43 (.I(rdata[4]),
    .Z(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input44 (.I(rdata[5]),
    .Z(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input45 (.I(rdata[6]),
    .Z(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(rdata[7]),
    .Z(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(rdata[8]),
    .Z(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(rdata[9]),
    .Z(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input49 (.I(reset),
    .Z(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(inst[13]),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(inst[14]),
    .Z(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input7 (.I(inst[15]),
    .Z(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(inst[1]),
    .Z(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(inst[2]),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net137),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I (.I(microcode),
    .ZN(microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q (.D(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .CLK(clknet_2_3__leaf_clk),
    .Q(microcode),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN),
    .A2(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .B(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_B),
    .C(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .ZN(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_147 (.ZN(net147),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_148 (.ZN(net148),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_149 (.ZN(net149),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_150 (.ZN(net150),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_151 (.ZN(net151),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_152 (.ZN(net152),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_153 (.ZN(net153),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_154 (.ZN(net154),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_155 (.ZN(net155),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_156 (.ZN(net156),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_157 (.ZN(net157),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_158 (.ZN(net158),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_159 (.ZN(net159),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_160 (.ZN(net160),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_161 (.ZN(net161),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_162 (.ZN(net162),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_163 (.ZN(net163),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_164 (.ZN(net164),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_165 (.ZN(net165),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_166 (.ZN(net166),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_167 (.ZN(net167),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_168 (.ZN(net168),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_169 (.ZN(net169),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_170 (.ZN(net170),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_171 (.ZN(net171),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_172 (.ZN(net172),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_173 (.ZN(net173),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_174 (.ZN(net174),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_175 (.ZN(net175),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_176 (.ZN(net176),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_177 (.ZN(net177),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_178 (.ZN(net178),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel minimax_179 (.ZN(net179),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .Z(op16_lw),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .ZN(op16_lw_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 op16_lwsp_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2 (.A1(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .A2(op16_lwsp),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D (.D(op16_slli_setrd),
    .CLK(clknet_2_3__leaf_clk),
    .Q(dly16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .ZN(op16_slli_setrd),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(net4),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2 (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2),
    .A3(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3),
    .A4(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B),
    .C(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A3),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A4(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A2_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_A2),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_A4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3 (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .A3(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN),
    .Z(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__and2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN),
    .ZN(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .A2(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .C(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A2),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .ZN(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .B1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .B2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand4_1_ZN_A3 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .ZN(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_A1),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__or2_2_Z (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .A2(net7),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .B1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or2_1_Z_A1),
    .B2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2 (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1),
    .Z(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_2_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B),
    .C(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_C),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z (.A1(net135),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN (.A1(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .A3(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_C_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(\pc_execute[8] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_C),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_A2),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__mux2_2_Z (.I0(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .I1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ),
    .S(\pc_execute[6] ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_B),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2 (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D (.D(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2 (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_A2),
    .B1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1),
    .B2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A2(\pc_execute[5] ),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_B1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .Z(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .A2(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN (.I(net10),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1 (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1),
    .A2(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .ZN(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .Z(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(net9),
    .Z(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D (.D(op16_slli_setrs),
    .CLK(clknet_2_3__leaf_clk),
    .Q(dly16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1),
    .A2(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .ZN(op16_slli_setrs),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .ZN(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN (.I(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .ZN(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1 (.A1(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2),
    .A2(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .ZN(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z (.I(dly16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_4_B_A1),
    .Z(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I (.I(op16_slli_setrs_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .Z(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output100 (.I(net100),
    .Z(aluX[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output101 (.I(net101),
    .Z(aluX[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output102 (.I(net102),
    .Z(aluX[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output103 (.I(net103),
    .Z(aluX[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output104 (.I(net104),
    .Z(aluX[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output105 (.I(net105),
    .Z(aluX[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output106 (.I(net106),
    .Z(aluX[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output107 (.I(net107),
    .Z(aluX[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output108 (.I(net108),
    .Z(aluX[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output109 (.I(net109),
    .Z(aluX[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output110 (.I(net110),
    .Z(aluX[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output111 (.I(net111),
    .Z(aluX[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output112 (.I(net112),
    .Z(aluX[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output113 (.I(net113),
    .Z(aluX[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output114 (.I(net114),
    .Z(aluX[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output115 (.I(net115),
    .Z(aluX[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output116 (.I(net116),
    .Z(aluX[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output117 (.I(net117),
    .Z(aluX[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output118 (.I(net118),
    .Z(aluX[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output119 (.I(net119),
    .Z(aluX[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output120 (.I(net120),
    .Z(aluX[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output121 (.I(net121),
    .Z(aluX[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output122 (.I(net122),
    .Z(aluX[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output123 (.I(net123),
    .Z(aluX[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output124 (.I(net124),
    .Z(aluX[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output125 (.I(net125),
    .Z(aluX[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output126 (.I(net126),
    .Z(inst_addr[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output127 (.I(net127),
    .Z(inst_addr[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output128 (.I(net128),
    .Z(inst_addr[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output129 (.I(net129),
    .Z(inst_addr[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output130 (.I(net130),
    .Z(inst_addr[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output131 (.I(net131),
    .Z(inst_addr[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output132 (.I(net132),
    .Z(inst_addr[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output133 (.I(net133),
    .Z(inst_addr[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output134 (.I(net134),
    .Z(inst_addr[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output135 (.I(net135),
    .Z(inst_addr[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output136 (.I(net136),
    .Z(inst_addr[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output137 (.I(net137),
    .Z(inst_regce),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output138 (.I(net138),
    .Z(rreq),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output139 (.I(net139),
    .Z(wb),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output140 (.I(net140),
    .Z(wmask[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output141 (.I(net141),
    .Z(wmask[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output142 (.I(net142),
    .Z(wmask[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output143 (.I(net143),
    .Z(wmask[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(addrD[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(addrD[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(addrD[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(addrD[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(addrD[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(addrD[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(addrS[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(addrS[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(addrS[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(addrS[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(addrS[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(addrS[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(addr[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(addr[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(addr[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(addr[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(addr[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(addr[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(addr[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(addr[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(addr[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(addr[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(addr[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(addr[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(addr[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(addr[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(addr[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(addr[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(addr[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(addr[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output80 (.I(net80),
    .Z(addr[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output81 (.I(net81),
    .Z(addr[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output82 (.I(net82),
    .Z(addr[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(addr[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output84 (.I(net84),
    .Z(addr[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output85 (.I(net85),
    .Z(addr[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output86 (.I(net86),
    .Z(addr[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output87 (.I(net87),
    .Z(addr[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output88 (.I(net88),
    .Z(addr[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output89 (.I(net89),
    .Z(addr[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output90 (.I(net90),
    .Z(addr[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output91 (.I(net91),
    .Z(addr[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output92 (.I(net92),
    .Z(addr[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output93 (.I(net93),
    .Z(addr[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output94 (.I(net94),
    .Z(aluX[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output95 (.I(net95),
    .Z(aluX[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output96 (.I(net96),
    .Z(aluX[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output97 (.I(net97),
    .Z(aluX[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output98 (.I(net98),
    .Z(aluX[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output99 (.I(net99),
    .Z(aluX[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I  (.I(\pc_execute[10] ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_execute[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .A2(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .B(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .B(\pc_execute[10] ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .A3(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S  (.I0(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .I1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .S(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN  (.A1(\pc_execute[8] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .C(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\pc_execute[9] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .B1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .B2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .B(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN  (.A1(\pc_execute[8] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B ),
    .C(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z),
    .A3(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .B(\pc_execute[8] ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S  (.I0(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .I1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .S(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net136),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN  (.A1(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .B1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .B2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .A3(net16),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_ZN_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(net126),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S  (.I0(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .I1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .S(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 \pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .A3(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ),
    .A4(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_execute[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_execute[11] ),
    .I1(\pc_fetch_dly[11] ),
    .S(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2  (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .A2(\pc_execute[11] ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .Z(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net4),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A4  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A4(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_A1 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1  (.A1(net127),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .B1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .B2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .ZN(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2  (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z ),
    .I1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .S(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I  (.I(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2  (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .ZN(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_execute[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_execute[1] ),
    .I1(\pc_fetch_dly[1] ),
    .S(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\pc_execute[1] ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net10),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .A2(\pc_execute[2] ),
    .A3(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_B2 ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ),
    .B(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .ZN(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(net16),
    .A2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A2 ),
    .B1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .B2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_B_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z ),
    .B(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\pc_execute[1] ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .B1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .B2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z  (.A1(net128),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I  (.I(\pc_execute[3] ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .C(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A1 ),
    .A2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3_ZN ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_C ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(net131),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A2 ),
    .B1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .B2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\pc_execute[4] ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2  (.A1(\pc_execute[4] ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN ),
    .B(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A1  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_execute[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN ),
    .A2(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .B(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .B(\pc_execute[3] ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .A4(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_A1),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A3(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A4(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net6),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z  (.I(net5),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ),
    .B1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1 ),
    .B2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .C(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C ),
    .ZN(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__and4_2_A3_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nor3_2_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_2_ZN_A1),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1 ),
    .B(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__oai22_1_ZN_A2),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai31_1_ZN  (.A1(net8),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_A1 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A2 ),
    .B(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A2_C ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A3  (.A1(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A2_A1),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A2_ZN),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ),
    .ZN(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .A3(net14),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net12),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A4(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .A4(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A4 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2  (.A1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_Z ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN ),
    .B1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1 ),
    .B2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2 ),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .A2(\pc_execute[4] ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(net131),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .Z(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A4_ZN ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_A2_ZN ),
    .B(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A3 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN ),
    .B1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_B_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .B2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .A2(\pc_execute[5] ),
    .A3(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .A3(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_2_A1_ZN),
    .B1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1 ),
    .B2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN  (.A1(\pc_execute[6] ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .B(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1 ),
    .C(\pc_execute[5] ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[6] ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_B2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai32_4_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2  (.A1(op16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A1_ZN),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi221_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xnor2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A2_ZN ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_Z ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1  (.A1(\pc_execute[3] ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A2(\pc_execute[2] ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .A2(\pc_execute[2] ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(net11),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand4_2_ZN_A2 ),
    .A3(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A4_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A4(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__nor4_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and3_1_Z_A3 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z ),
    .B(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z  (.A1(net130),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ),
    .Z(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3  (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ),
    .A3(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN ),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .A2(microcode_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__aoi211_2_ZN_A2),
    .ZN(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_ZN ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\pc_execute[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_execute[7] ),
    .I1(\pc_fetch_dly[7] ),
    .S(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_2_Z  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(net13),
    .A2(\pc_execute[7] ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2  (.A1(net13),
    .A2(\pc_execute[7] ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .B1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1 ),
    .B2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(net134),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1 ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor2_2_A1  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .Z(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_A2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_A1 ),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A1 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_A2 ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S  (.I0(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .I1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .S(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1_gf180mcu_fd_sc_mcu7t5v0__nor2_1_ZN  (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A2 ),
    .ZN(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_I1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I  (.I(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z ),
    .Z(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__mux2_2_S_Z_gf180mcu_fd_sc_mcu7t5v0__buf_4_I_Z ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net135),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \pc_execute[8]_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I  (.I(\pc_execute[8] ),
    .ZN(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1  (.A1(\pc_execute[9] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .B(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_B ),
    .ZN(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_1  (.A1(\pc_execute[9] ),
    .A2(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .B(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_ZN_B_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_ZN_C ),
    .ZN(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B  (.A1(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B2 ),
    .A2(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .B(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN ),
    .ZN(\pc_execute[10]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__nor3_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z  (.A1(net136),
    .A2(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_2_A2_B1_gf180mcu_fd_sc_mcu7t5v0__and2_1_Z_A2 ),
    .Z(\pc_execute[9]_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_B_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\pc_fetch_dly[10] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .B1(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net18),
    .ZN(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(net41),
    .A2(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .ZN(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .A2(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .ZN(net118),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2  (.A1(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ),
    .A2(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net95),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(net63),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .ZN(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_fetch_dly[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[10] ),
    .I1(net126),
    .S(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_fetch_dly[10] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .ZN(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\pc_fetch_dly[11] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .B1(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net19),
    .ZN(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2  (.A1(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A2_A1 ),
    .A2(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net96),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_fetch_dly[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[11] ),
    .I1(net127),
    .S(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[11]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_fetch_dly[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .A2(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(net128),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .ZN(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2  (.A1(net129),
    .A2(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .Z(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A3  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_B2 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A1_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor3_2_A3_A2 ),
    .A3(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z ),
    .ZN(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_Z_gf180mcu_fd_sc_mcu7t5v0__aoi21_1_A2_B ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_fetch_dly[1] ),
    .A2(net138),
    .ZN(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1  (.A1(\pc_fetch_dly[1] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .ZN(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ),
    .A2(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ),
    .ZN(net105),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(net73),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B1(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net28),
    .ZN(\pc_fetch_dly[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1  (.A1(\pc_fetch_dly[2] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .B1(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B2(net84),
    .C1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .C2(net39),
    .ZN(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(net69),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .ZN(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ),
    .ZN(net101),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(net24),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z),
    .ZN(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_3_I  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .ZN(net116),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\pc_fetch_dly[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[2] ),
    .I1(net129),
    .S(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1  (.I0(\pc_execute[2] ),
    .I1(\pc_fetch_dly[2] ),
    .S(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .Z(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_execute[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\pc_fetch_dly[3] ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net42),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .Z(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net119),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_A1 ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .B1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .B2(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_A1 ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_B ),
    .A2(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi211_1_A2_C_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .ZN(net87),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_fetch_dly[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .A2(net138),
    .B(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net130),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1  (.A1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .A2(\pc_execute[3]_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_2_A3_A1 ),
    .A3(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ),
    .Z(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(net128),
    .A2(net129),
    .A3(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_A1_gf180mcu_fd_sc_mcu7t5v0__xor2_1_Z_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3_gf180mcu_fd_sc_mcu7t5v0__inv_1_ZN  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A1_A3_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_fetch_dly[3] ),
    .A2(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1  (.A1(\pc_fetch_dly[3] ),
    .A2(net138),
    .ZN(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\pc_fetch_dly[4] ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net43),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net120),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .B1(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .B2(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C2 ),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ),
    .A2(\dra[2]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1_gf180mcu_fd_sc_mcu7t5v0__oai221_4_A1_B1 ),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_A2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .ZN(net88),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_fetch_dly[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN  (.A1(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .A2(net138),
    .B(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_ZN  (.I(net131),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__oai21_1_ZN_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1  (.I0(\pc_execute[4] ),
    .I1(\pc_fetch_dly[4] ),
    .S(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .Z(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\pc_execute[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_fetch_dly[4] ),
    .A2(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .ZN(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1  (.A1(\pc_fetch_dly[5] ),
    .A2(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .B1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .B2(net44),
    .ZN(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B  (.A1(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A2 ),
    .B(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN ),
    .ZN(net121),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN  (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B2 ),
    .A2(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_A1_A2),
    .B1(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .B2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .ZN(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN  (.A1(\dra[1]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand3_1_ZN_A2 ),
    .A2(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__xor3_1_A3_A1_gf180mcu_fd_sc_mcu7t5v0__oai21_2_A1_A2 ),
    .A3(bubble1_gf180mcu_fd_sc_mcu7t5v0__or3_2_A2_Z_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_1_A1_ZN),
    .ZN(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_ZN_B1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1_gf180mcu_fd_sc_mcu7t5v0__inv_1_I  (.I(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_2_B_A1 ),
    .ZN(net89),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\pc_fetch_dly[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[5] ),
    .I1(net132),
    .S(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1  (.I0(\pc_execute[5] ),
    .I1(\pc_fetch_dly[5] ),
    .S(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .Z(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[5]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\pc_execute[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1  (.A1(\pc_fetch_dly[6] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_A2 ),
    .B1(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B2(net90),
    .C1(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .C2(net45),
    .ZN(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I  (.I(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .ZN(net122),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\pc_fetch_dly[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[6] ),
    .I1(net133),
    .S(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1  (.I0(\pc_execute[6] ),
    .I1(\pc_fetch_dly[6] ),
    .S(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .Z(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[6]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\pc_execute[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1  (.A1(\pc_fetch_dly[7] ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B2(net91),
    .C1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .C2(net46),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(net68),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1  (.A1(net67),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .ZN(net99),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2  (.A1(net66),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .ZN(net98),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3  (.A1(net65),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .ZN(net97),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4  (.A1(net62),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .ZN(net94),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_3_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .ZN(net100),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2  (.A1(net70),
    .A2(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .ZN(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .ZN(net112),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .ZN(net111),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .ZN(net110),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .ZN(net109),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_4  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_1_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .ZN(net108),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_1_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_4_ZN),
    .ZN(net107),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .ZN(net106),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .ZN(net104),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .ZN(net103),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_4  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_2_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_2_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .ZN(net102),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN),
    .ZN(net117),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_1  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_1_ZN),
    .ZN(net115),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_2  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_2_ZN),
    .ZN(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_2_A1_3  (.A1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_ZN_gf180mcu_fd_sc_mcu7t5v0__buf_2_I_Z ),
    .A2(dly16_lw_gf180mcu_fd_sc_mcu7t5v0__or2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A2_3_ZN),
    .ZN(net113),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .ZN(net123),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\pc_fetch_dly[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[7] ),
    .I1(net134),
    .S(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1  (.A1(\pc_fetch_dly[8] ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B2(net92),
    .C1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .C2(net47),
    .ZN(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I  (.I(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_A1_ZN ),
    .ZN(net124),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\pc_fetch_dly[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[8] ),
    .I1(net135),
    .S(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1  (.A1(\pc_fetch_dly[8] ),
    .A2(\pc_fetch_dly[2]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .ZN(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B  (.A1(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_A1 ),
    .A2(inst_regce_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D),
    .B(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN ),
    .ZN(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[8]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__oai21_1_B_ZN ),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\pc_execute[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1  (.A1(\pc_fetch_dly[9] ),
    .A2(\pc_fetch_dly[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_A2 ),
    .B1(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_B1 ),
    .B2(net93),
    .C1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__or2_1_A1_A2),
    .C2(net48),
    .ZN(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__inv_2_I  (.I(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__aoi222_2_A1_ZN ),
    .ZN(net125),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q  (.D(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_fetch_dly[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z  (.I(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .Z(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__dffq_1_Q_D ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0  (.I0(\pc_fetch_dly[9] ),
    .I1(net136),
    .S(\pc_fetch_dly[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1  (.I0(\pc_execute[9] ),
    .I1(\pc_fetch_dly[9] ),
    .S(\pc_execute[7]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I0_S ),
    .Z(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I  (.I(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z ),
    .Z(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D  (.D(\pc_fetch_dly[9]_gf180mcu_fd_sc_mcu7t5v0__mux2_2_I1_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z ),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\pc_execute[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(net49),
    .Z(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__clkinv_1_I (.I(reset_gf180mcu_fd_sc_mcu7t5v0__buf_1_I_Z),
    .ZN(\pc_execute[11]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__and2_1_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I (.I(net49),
    .Z(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__buf_1_I (.I(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .Z(\pc_execute[1]_gf180mcu_fd_sc_mcu7t5v0__xor2_1_A2_Z_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B1_ZN_gf180mcu_fd_sc_mcu7t5v0__nor2_2_A2_A1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1 (.A1(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z),
    .A2(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_A2),
    .ZN(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_ZN),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_ZN_gf180mcu_fd_sc_mcu7t5v0__dffq_1_D (.D(reset_gf180mcu_fd_sc_mcu7t5v0__clkbuf_1_I_Z_gf180mcu_fd_sc_mcu7t5v0__nor2_4_A1_ZN),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net134),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rreq_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(\pc_fetch_dly[4]_gf180mcu_fd_sc_mcu7t5v0__nand2_1_A1_A2 ),
    .Z(net138),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .Z(net139),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z (.A1(\dra[0]_gf180mcu_fd_sc_mcu7t5v0__aoi221_1_A1_C ),
    .A2(\pc_fetch_dly[10]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_A1_B1 ),
    .A3(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3),
    .Z(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3_gf180mcu_fd_sc_mcu7t5v0__oai211_1_ZN (.A1(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A1),
    .A2(dly16_slli_setrd_gf180mcu_fd_sc_mcu7t5v0__nor3_1_A2_A3),
    .B(\dra[4]_gf180mcu_fd_sc_mcu7t5v0__aoi222_1_B2_C1_gf180mcu_fd_sc_mcu7t5v0__nand2_1_ZN_A1 ),
    .C(\dra[3]_gf180mcu_fd_sc_mcu7t5v0__aoi22_1_B2_ZN_gf180mcu_fd_sc_mcu7t5v0__nand4_1_A3_A2 ),
    .ZN(wb_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_I_gf180mcu_fd_sc_mcu7t5v0__or3_1_Z_A3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z (.I(net143),
    .Z(net142),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_1 (.I(net143),
    .Z(net140),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wmask_gf180mcu_fd_sc_mcu7t5v0__buf_1_Z_2 (.I(net143),
    .Z(net141),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign inst_addr[0] = net147;
 assign wdata[0] = net173;
 assign wdata[10] = net162;
 assign wdata[11] = net161;
 assign wdata[12] = net159;
 assign wdata[13] = net158;
 assign wdata[14] = net157;
 assign wdata[15] = net156;
 assign wdata[16] = net155;
 assign wdata[17] = net154;
 assign wdata[18] = net153;
 assign wdata[19] = net152;
 assign wdata[1] = net172;
 assign wdata[20] = net151;
 assign wdata[21] = net150;
 assign wdata[22] = net179;
 assign wdata[23] = net178;
 assign wdata[24] = net177;
 assign wdata[25] = net176;
 assign wdata[26] = net175;
 assign wdata[27] = net174;
 assign wdata[28] = net171;
 assign wdata[29] = net160;
 assign wdata[2] = net170;
 assign wdata[30] = net149;
 assign wdata[31] = net148;
 assign wdata[3] = net169;
 assign wdata[4] = net168;
 assign wdata[5] = net167;
 assign wdata[6] = net166;
 assign wdata[7] = net165;
 assign wdata[8] = net164;
 assign wdata[9] = net163;
endmodule
