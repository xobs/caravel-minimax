* NGSPICE file created from RAM32_1RW1R.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latq_1 D E Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_1 EN I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__icgtp_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__icgtp_1 CLK E TE Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

.subckt RAM32_1RW1R A0[0] A0[1] A0[2] A0[3] A0[4] A1[0] A1[1] A1[2] A1[3] A1[4] CLK
+ Di0[0] Di0[10] Di0[11] Di0[12] Di0[13] Di0[14] Di0[15] Di0[16] Di0[17] Di0[18] Di0[19]
+ Di0[1] Di0[20] Di0[21] Di0[22] Di0[23] Di0[24] Di0[25] Di0[26] Di0[27] Di0[28] Di0[29]
+ Di0[2] Di0[30] Di0[31] Di0[3] Di0[4] Di0[5] Di0[6] Di0[7] Di0[8] Di0[9] Do0[0] Do0[10]
+ Do0[11] Do0[12] Do0[13] Do0[14] Do0[15] Do0[16] Do0[17] Do0[18] Do0[19] Do0[1] Do0[20]
+ Do0[21] Do0[22] Do0[23] Do0[24] Do0[25] Do0[26] Do0[27] Do0[28] Do0[29] Do0[2] Do0[30]
+ Do0[31] Do0[3] Do0[4] Do0[5] Do0[6] Do0[7] Do0[8] Do0[9] Do1[0] Do1[10] Do1[11]
+ Do1[12] Do1[13] Do1[14] Do1[15] Do1[16] Do1[17] Do1[18] Do1[19] Do1[1] Do1[20] Do1[21]
+ Do1[22] Do1[23] Do1[24] Do1[25] Do1[26] Do1[27] Do1[28] Do1[29] Do1[2] Do1[30] Do1[31]
+ Do1[3] Do1[4] Do1[5] Do1[6] Do1[7] Do1[8] Do1[9] EN0 EN1 VDD VSS WE0[0] WE0[1] WE0[2]
+ WE0[3]
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_552 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_541 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_530 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_596 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_585 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_574 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_563 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.DEC1.AND0 SLICE\[2\].RAM8.DEC1.A_buf\[0\] SLICE\[2\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC1.A_buf\[2\] SLICE\[2\].RAM8.DEC1.EN_buf_N SLICE\[2\].RAM8.WORD\[0\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XSLICE\[0\].RAM8.DEC1.ENBUF SLICE\[0\].RAM8.DEC1.EN SLICE\[0\].RAM8.DEC1.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_29_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_10_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_28_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_19_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_33_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[2\].W.SEL0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_6_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_6_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BYTE\[1\].FLOATBUF1\[11\].Z Do1_REG.CLKBUF\[1\]
+ Do1[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_16_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_32_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_22_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_30_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BYTE\[3\].FLOATBUF0\[30\].Z Do0_REG.CLKBUF\[3\]
+ Do0[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_30_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC0.INV3 SLICE\[3\].RAM8.DEC0.A_buf\[1\] SLICE\[3\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\].X SLICE\[3\].RAM8.DEC1.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_21_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_8_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_12_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_33_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_12_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[0\].W.SEL1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.AND4 SLICE\[1\].RAM8.DEC0.A_buf_N\[0\] SLICE\[1\].RAM8.DEC0.A_buf_N\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[4\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[27\].__cell__ BYTE\[3\].FLOATBUF0\[27\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[27\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[0\].FLOATBUF1\[5\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[5\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_701 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_745 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_734 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_723 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_712 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_778 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_767 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_756 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_33_789 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_9_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_9_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_5_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_24_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[3\].FLOATBUF1\[24\].__cell__ BYTE\[3\].FLOATBUF1\[24\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[24\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_520 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_553 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_542 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_531 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_33_586 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_575 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_564 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_597 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_20_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_15_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_9_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_5_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.AND1 zero_ SLICE\[2\].RAM8.DEC1.A_buf_N\[1\] SLICE\[2\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[1\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_19_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_19_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_1_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[1\].W.SEL0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_2_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF0\[0\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[0\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_22_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BYTE\[0\].FLOATBUF0\[3\].Z Do0_REG.CLKBUF\[0\]
+ Do0[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_21_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_18_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[24\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[24\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_25_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.ENBUF SLICE\[0\].RAM8.DEC0.EN SLICE\[0\].RAM8.DEC0.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BYTE\[2\].FLOATBUF1\[23\].Z Do1_REG.CLKBUF\[2\]
+ Do1[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_20_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_0_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_469 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_458 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_29_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.INV4 SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.DEC0.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtap_8_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_11_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[24\].__cell__ Di0[24] DIBUF\[24\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_12_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[31\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[31\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_33_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_12_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.AND5 SLICE\[1\].RAM8.DEC0.A_buf_N\[1\] SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[5\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XBYTE\[2\].FLOATBUF0\[19\].__cell__ BYTE\[2\].FLOATBUF0\[19\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[19\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_702 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[7\].W.SEL1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_735 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_724 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_713 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_768 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_757 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_746 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_779 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_0_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BYTE\[3\].FLOATBUF1\[24\].Z Do1_REG.CLKBUF\[3\]
+ Do1[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_9_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_9_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDIBUF\[8\].__cell__ Di0[8] DIBUF\[8\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_24_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_24_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF0\[10\].__cell__ BYTE\[1\].FLOATBUF0\[10\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[10\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_510 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_543 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_532 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_521 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[0\].W.SEL0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_33_587 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_576 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_565 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_554 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_598 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_20_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBYTE\[2\].FLOATBUF1\[16\].__cell__ BYTE\[2\].FLOATBUF1\[16\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[16\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_0_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_5_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.DEC1.AND2 zero_ SLICE\[2\].RAM8.DEC1.A_buf_N\[0\] SLICE\[2\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[2\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_29_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[10\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[10\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_2_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF0\[4\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[4\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[21\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[21\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_13_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BYTE\[1\].FLOATBUF0\[15\].Z Do0_REG.CLKBUF\[1\]
+ Do0[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_1_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_21_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[2\].FLOATBUF0\[17\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[17\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_18_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[28\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[28\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_7_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtap_11_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[14\].__cell__ Di0[14] DIBUF\[14\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_16_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_22_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_9_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_29_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[6\].W.SEL1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_8_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_11_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_27_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_31_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.CLKBUF.__cell__ CLKBUF.X SLICE\[2\].RAM8.CLKBUF.X VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_31_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.AND6 SLICE\[1\].RAM8.DEC0.A_buf_N\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[6\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_0_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BYTE\[2\].FLOATBUF0\[16\].Z Do0_REG.CLKBUF\[2\]
+ Do0[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_26_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_21_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_17_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtap_13_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_736 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_725 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_714 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_703 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_769 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_758 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_747 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_32_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_24_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_24_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_511 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_500 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_544 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_533 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_577 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_566 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_555 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF1\[3\].__cell__ BYTE\[0\].FLOATBUF1\[3\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[3\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_599 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_588 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_20_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_8_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_9_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_5_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.DEC1.AND3 zero_ SLICE\[2\].RAM8.DEC1.A_buf\[1\] SLICE\[2\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[3\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_29_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A SLICE\[3\].RAM8.WEBUF\[2\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_1_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_6_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[14\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[14\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[7\].__cell__ BYTE\[0\].FLOATBUF0\[7\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[7\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_19_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_19_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtap_11_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[5\].W.SEL1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_31_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_16_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_32_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_13_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_9_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BYTE\[1\].FLOATBUF1\[9\].Z Do1_REG.CLKBUF\[1\]
+ Do1[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_29_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_15_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_15_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BYTE\[3\].FLOATBUF0\[28\].Z Do0_REG.CLKBUF\[3\]
+ Do0[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[1\].RAM8.DEC0.AND7 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[7\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_0_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\].X SLICE\[3\].RAM8.DEC1.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_26_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_26_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_17_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_17_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_33_726 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_715 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_704 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_759 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_748 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_737 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_24_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_0_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_0_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_26_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.CLKBUF.__cell__ CLKBUF.X SLICE\[0\].RAM8.CLKBUF.X VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_24_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_501 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_534 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_523 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_512 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[26\].__cell__ BYTE\[3\].FLOATBUF0\[26\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[26\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_578 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_567 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_556 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_545 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_589 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_20_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_14_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_9_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.AND4 SLICE\[2\].RAM8.DEC1.A_buf_N\[0\] SLICE\[2\].RAM8.DEC1.A_buf_N\[1\]
+ SLICE\[2\].RAM8.DEC1.A_buf\[2\] SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[4\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_10_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_19_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_1_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_13_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[4\].W.SEL1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_28_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_1_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_18_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_25_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_32_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BYTE\[0\].FLOATBUF0\[1\].Z Do0_REG.CLKBUF\[0\]
+ Do0[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_22_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_20_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_13_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BYTE\[2\].FLOATBUF1\[21\].Z Do1_REG.CLKBUF\[2\]
+ Do1[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_3_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_15_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_0_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_26_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_727 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_716 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_705 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_749 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_738 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_32_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_9_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_23_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDIBUF\[23\].__cell__ Di0[23] DIBUF\[23\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\].X SLICE\[0\].RAM8.DEC1.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_8_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_4_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_24_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_502 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_33_535 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_524 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_568 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_557 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_546 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_579 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[2\].FLOATBUF0\[18\].__cell__ BYTE\[2\].FLOATBUF0\[18\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[18\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[3\].W.SEL1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_0_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_14_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.AND5 SLICE\[2\].RAM8.DEC1.A_buf_N\[1\] SLICE\[2\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC1.A_buf\[2\] SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[5\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_19_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDIBUF\[7\].__cell__ Di0[7] DIBUF\[7\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_33_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_6_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_1_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_27_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.ENBUF SLICE\[3\].RAM8.DEC1.EN SLICE\[3\].RAM8.DEC1.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XWEBUF\[3\].__cell__ WE0[3] SLICE\[0\].RAM8.WEBUF\[3\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_25_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_24_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BYTE\[1\].FLOATBUF0\[13\].Z Do0_REG.CLKBUF\[1\]
+ Do0[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_16_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_30_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC0.INV1 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_21_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_27_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[13\].__cell__ Di0[13] DIBUF\[13\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_0_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_26_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_717 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_706 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_739 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_728 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_32_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[2\].W.SEL1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_26_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_9_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_9_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[25\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[25\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_14_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_8_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_24_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_525 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_514 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_503 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_569 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_558 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_547 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_536 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.AND6 SLICE\[2\].RAM8.DEC1.A_buf_N\[0\] SLICE\[2\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC1.A_buf\[2\] SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[6\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_29_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_19_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_23_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_25_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_6_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XBYTE\[0\].FLOATBUF1\[2\].__cell__ BYTE\[0\].FLOATBUF1\[2\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[2\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_27_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BYTE\[0\].FLOATBUF1\[6\].Z Do1_REG.CLKBUF\[0\]
+ Do1[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_18_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_11_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A SLICE\[3\].RAM8.WEBUF\[1\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_25_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF0\[6\].__cell__ BYTE\[0\].FLOATBUF0\[6\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[6\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_18_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_30_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC0.INV2 SLICE\[1\].RAM8.DEC0.A_buf\[1\] SLICE\[1\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_10_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_10_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_10_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_29_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.ENBUF SLICE\[3\].RAM8.DEC0.EN SLICE\[3\].RAM8.DEC0.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A SLICE\[2\].RAM8.WEBUF\[3\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_12_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[1\].W.SEL1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_33_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X SLICE\[1\].RAM8.DEC0.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_21_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[22\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[22\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_718 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_707 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_729 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_9_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BYTE\[3\].FLOATBUF0\[26\].Z Do0_REG.CLKBUF\[3\]
+ Do0[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_29_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[29\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[29\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_526 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_515 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_559 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_548 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_537 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_22_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_8_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_30_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.DEC1.AND7 SLICE\[2\].RAM8.DEC1.A_buf\[0\] SLICE\[2\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC1.A_buf\[2\] SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.WORD\[7\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.AND0 SLICE\[0\].RAM8.DEC1.A_buf\[0\] SLICE\[0\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC1.A_buf\[2\] SLICE\[0\].RAM8.DEC1.EN_buf_N SLICE\[0\].RAM8.WORD\[0\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_4_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_6_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_20_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[25\].__cell__ BYTE\[3\].FLOATBUF0\[25\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[25\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_27_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XA0BUF\[4\].__cell__ A0[4] A0BUF\[4\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF1\[12\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[12\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_11_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[1\].RAM8.WORD\[0\].W.SEL1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[2\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\].X SLICE\[2\].RAM8.DEC1.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[19\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[19\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.DEC0.INV3 SLICE\[1\].RAM8.DEC0.A_buf\[1\] SLICE\[1\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo1_REG.Do_CLKBUF\[3\] Do1_REG.CLK_buf Do1_REG.CLKBUF\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_10_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_19_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_33_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_26_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BYTE\[2\].FLOATBUF1\[19\].Z Do1_REG.CLKBUF\[2\]
+ Do1[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_21_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_708 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_719 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_32_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_0_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_31_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_29_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_28_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_8_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_33_516 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_505 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_549 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_538 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_527 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_7_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_8_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_30_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.AND1 zero_ SLICE\[0\].RAM8.DEC1.A_buf_N\[1\] SLICE\[0\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[1\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[22\].__cell__ Di0[22] DIBUF\[22\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_33_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_6_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_25_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_1_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_27_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[17\].__cell__ BYTE\[2\].FLOATBUF0\[17\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[17\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_11_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[6\].__cell__ Di0[6] DIBUF\[6\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_6_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_15_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[0\].FLOATBUF1\[0\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[0\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_22_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.DEC0.INV4 SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.DEC0.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_10_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[7\].W.SEL1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_10_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XWEBUF\[2\].__cell__ WE0[2] SLICE\[0\].RAM8.WEBUF\[2\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_12_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_7_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[3\] BYTE\[1\].FLOATBUF0\[11\].Z Do0_REG.CLKBUF\[1\]
+ Do0[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_7_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_23_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BYTE\[3\].FLOATBUF1\[31\].Z Do1_REG.CLKBUF\[3\]
+ Do1[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_33_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[1\].FLOATBUF1\[9\].__cell__ BYTE\[1\].FLOATBUF1\[9\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[9\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_709 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_0_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_31_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtap_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.INV1 SLICE\[2\].RAM8.DEC1.A_buf\[0\] SLICE\[2\].RAM8.DEC1.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDIBUF\[12\].__cell__ Di0[12] DIBUF\[12\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_33_517 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_539 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_528 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_7_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.AND2 zero_ SLICE\[0\].RAM8.DEC1.A_buf_N\[0\] SLICE\[0\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[2\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_390 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_33_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_13_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_1_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X SLICE\[3\].RAM8.DEC0.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_18_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[6\].W.SEL1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_18_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_30_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BYTE\[0\].FLOATBUF1\[4\].Z Do1_REG.CLKBUF\[0\]
+ Do1[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_29_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[0\].FLOATBUF1\[1\].__cell__ BYTE\[0\].FLOATBUF1\[1\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[1\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF1\[4\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[4\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_21_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_10_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_10_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_29_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[7\] BYTE\[2\].FLOATBUF0\[23\].Z Do0_REG.CLKBUF\[2\]
+ Do0[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_12_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_12_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_23_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A SLICE\[3\].RAM8.WEBUF\[0\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_11_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[5\].__cell__ BYTE\[0\].FLOATBUF0\[5\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[5\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_9_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_29_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A SLICE\[2\].RAM8.WEBUF\[2\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC1.INV2 SLICE\[2\].RAM8.DEC1.A_buf\[1\] SLICE\[2\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_4_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_529 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_518 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[3\].FLOATBUF1\[31\].__cell__ BYTE\[3\].FLOATBUF1\[31\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[31\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_15_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_14_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[0\] BYTE\[3\].FLOATBUF0\[24\].Z Do0_REG.CLKBUF\[3\]
+ Do0[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_34_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_27_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_27_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.AND3 zero_ SLICE\[0\].RAM8.DEC1.A_buf\[1\] SLICE\[0\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[3\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_10_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_315 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[5\].W.SEL1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_19_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_27_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XBYTE\[3\].FLOATBUF0\[30\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[30\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_690 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_3_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[3\].FLOATBUF0\[24\].__cell__ BYTE\[3\].FLOATBUF0\[24\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[24\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_3_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XA0BUF\[3\].__cell__ A0[3] A0BUF\[3\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_7_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDIBUF\[31\].__cell__ Di0[31] DIBUF\[31\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\].X SLICE\[2\].RAM8.DEC1.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_33_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.Do_CLKBUF\[1\] Do1_REG.CLK_buf Do1_REG.CLKBUF\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_21_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_9_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BYTE\[2\].FLOATBUF1\[17\].Z Do1_REG.CLKBUF\[2\]
+ Do1[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.DEC1.INV3 SLICE\[2\].RAM8.DEC1.A_buf\[1\] SLICE\[2\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[3\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[3\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_519 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[20\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[20\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[4\].W.SEL1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_7_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[2\].FLOATBUF1\[23\].__cell__ BYTE\[2\].FLOATBUF1\[23\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[23\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_30_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF0\[16\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[16\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC1.AND4 SLICE\[0\].RAM8.DEC1.A_buf_N\[0\] SLICE\[0\].RAM8.DEC1.A_buf_N\[1\]
+ SLICE\[0\].RAM8.DEC1.A_buf\[2\] SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[4\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_10_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[27\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[27\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_4_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_4_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_6_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_20_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_13_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND0 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf_N SLICE\[2\].RAM8.WORD\[0\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xtap_6_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_13_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_27_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_18_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_11_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_4_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_680 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_691 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDIBUF\[21\].__cell__ Di0[21] DIBUF\[21\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_32_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_3_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XTIE1\[3\].__cell__ BYTE\[3\].FLOATBUF1\[24\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_22_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[16\].__cell__ BYTE\[2\].FLOATBUF0\[16\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[16\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_29_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_23_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_17_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[5\].__cell__ Di0[5] DIBUF\[5\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xtap_33_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_17_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[3\].W.SEL1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[1\] BYTE\[1\].FLOATBUF0\[9\].Z Do0_REG.CLKBUF\[1\]
+ Do0[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_0_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_16_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_31_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BYTE\[3\].FLOATBUF1\[29\].Z Do1_REG.CLKBUF\[3\]
+ Do1[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XWEBUF\[1\].__cell__ WE0[1] SLICE\[0\].RAM8.WEBUF\[1\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_16_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC1.INV4 SLICE\[2\].RAM8.DEC1.EN_buf SLICE\[2\].RAM8.DEC1.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XBYTE\[1\].FLOATBUF0\[13\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[13\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_509 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[7\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[7\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_7_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[8\].__cell__ BYTE\[1\].FLOATBUF1\[8\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[8\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_14_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[7\].W.SEL0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_30_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF1\[15\].__cell__ BYTE\[1\].FLOATBUF1\[15\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[15\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC1.AND5 SLICE\[0\].RAM8.DEC1.A_buf_N\[1\] SLICE\[0\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC1.A_buf\[2\] SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[5\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_382 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_371 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_360 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_393 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_3_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND1 zero_ SLICE\[2\].RAM8.DEC0.A_buf_N\[1\] SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[1\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_6_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_13_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_32_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[11\].__cell__ Di0[11] DIBUF\[11\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_11_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_24_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_681 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_670 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_692 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_32_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X SLICE\[3\].RAM8.DEC0.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_15_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_3_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_3_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFBUFENBUF1\[3\].__cell__ EN1 BYTE\[3\].FLOATBUF1\[24\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_22_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[2\].W.SEL1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_12_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_7_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_16_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.Do_CLKBUF\[3\] Do0_REG.CLK_buf Do0_REG.CLKBUF\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BYTE\[0\].FLOATBUF1\[2\].Z Do1_REG.CLKBUF\[0\]
+ Do1[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_17_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[5\] BYTE\[2\].FLOATBUF0\[21\].Z Do0_REG.CLKBUF\[2\]
+ Do0[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[0\].FLOATBUF1\[0\].__cell__ BYTE\[0\].FLOATBUF1\[0\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[0\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtap_9_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_9_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_14_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[6\].W.SEL0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_16_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_31_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_520 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_4_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_7_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF0\[4\].__cell__ BYTE\[0\].FLOATBUF0\[4\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[4\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_14_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_30_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_30_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_34_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_27_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_27_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC1.AND0 A1BUF\[3\].X A1BUF\[4\].X DEC1.EN_N SLICE\[0\].RAM8.DEC1.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
XSLICE\[0\].RAM8.DEC1.AND6 SLICE\[0\].RAM8.DEC1.A_buf_N\[0\] SLICE\[0\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC1.A_buf\[2\] SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[6\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_4_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_350 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_383 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_372 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_361 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_394 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A SLICE\[2\].RAM8.WEBUF\[1\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_6_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_13_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND2 zero_ SLICE\[2\].RAM8.DEC0.A_buf_N\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[2\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_6_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_32_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[3\].FLOATBUF1\[30\].__cell__ BYTE\[3\].FLOATBUF1\[30\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[30\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_0_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_11_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A SLICE\[1\].RAM8.WEBUF\[3\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_4_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[1\].W.SEL1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_7_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_671 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_660 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_693 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_682 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_30_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_23_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_12_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BYTE\[1\].FLOATBUF1\[14\].Z Do1_REG.CLKBUF\[1\]
+ Do1[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[5\].W.SEL0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X SLICE\[0\].RAM8.DEC0.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_4_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_25_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_9_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_14_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.ENBUF SLICE\[1\].RAM8.DEC1.EN SLICE\[1\].RAM8.DEC1.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_31_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XA0BUF\[2\].__cell__ A0[2] A0BUF\[2\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_16_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_32_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[30\].__cell__ Di0[30] DIBUF\[30\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_8_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_22_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_521 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_0_510 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_13_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_34_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_27_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_1_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC1.AND1 DEC1.A_N\[1\] A1BUF\[3\].X DEC1.EN SLICE\[1\].RAM8.DEC1.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XSLICE\[0\].RAM8.DEC1.AND7 SLICE\[0\].RAM8.DEC1.A_buf\[0\] SLICE\[0\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC1.A_buf\[2\] SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.WORD\[7\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_10_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_340 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_373 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_362 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_351 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_395 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_384 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_6_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND3 zero_ SLICE\[2\].RAM8.DEC0.A_buf\[1\] SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[3\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_6_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[0\].RAM8.WORD\[0\].W.SEL1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[2\].FLOATBUF1\[22\].__cell__ BYTE\[2\].FLOATBUF1\[22\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[22\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_1_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\].X SLICE\[1\].RAM8.DEC1.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XTIE_ZERO_zero_ zero_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xfill_24_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_661 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_650 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_694 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_683 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_672 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[4\].W.SEL0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_18_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_22_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[6\] BYTE\[0\].FLOATBUF0\[6\].Z Do0_REG.CLKBUF\[0\]
+ Do0[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.DEC1.AND0 SLICE\[3\].RAM8.DEC1.A_buf\[0\] SLICE\[3\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC1.A_buf\[2\] SLICE\[3\].RAM8.DEC1.EN_buf_N SLICE\[3\].RAM8.WORD\[0\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xfill_33_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_491 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[3\].FLOATBUF0\[24\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[24\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_11_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_17_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[20\].__cell__ Di0[20] DIBUF\[20\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_21_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_25_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XTIE1\[2\].__cell__ BYTE\[2\].FLOATBUF1\[16\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_21_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_9_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_14_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_29_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_28_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_522 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_0_511 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_500 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[4\].__cell__ Di0[4] DIBUF\[4\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_7_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_14_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_34_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_27_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BYTE\[3\].FLOATBUF1\[27\].Z Do1_REG.CLKBUF\[3\]
+ Do1[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_27_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDEC1.AND2 DEC1.A_N\[0\] A1BUF\[4\].X DEC1.EN SLICE\[2\].RAM8.DEC1.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
Xfill_4_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_4_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_341 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_330 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.ENBUF SLICE\[1\].RAM8.DEC0.EN SLICE\[1\].RAM8.DEC0.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_374 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_363 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_352 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_396 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_385 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_17_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XWEBUF\[0\].__cell__ WE0[0] SLICE\[0\].RAM8.WEBUF\[0\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND4 SLICE\[2\].RAM8.DEC0.A_buf_N\[0\] SLICE\[2\].RAM8.DEC0.A_buf_N\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[4\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_5_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_13_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[3\].W.SEL0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_1_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[14\].__cell__ BYTE\[1\].FLOATBUF1\[14\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[14\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_11_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_26_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_11_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_662 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_651 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_640 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_695 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_684 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_673 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_30_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[10\].__cell__ Di0[10] DIBUF\[10\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XBYTE\[2\].FLOATBUF0\[21\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[21\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.DEC1.AND1 zero_ SLICE\[3\].RAM8.DEC1.A_buf_N\[1\] SLICE\[3\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[1\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_12_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_470 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_20_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_25_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_11_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[28\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[28\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_17_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_21_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFBUFENBUF1\[2\].__cell__ EN1 BYTE\[2\].FLOATBUF1\[16\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_21_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.Do_CLKBUF\[1\] Do0_REG.CLK_buf Do0_REG.CLKBUF\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_16_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_31_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BYTE\[0\].FLOATBUF1\[0\].Z Do1_REG.CLKBUF\[0\]
+ Do1[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_29_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_22_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_512 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_501 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.INV1 SLICE\[0\].RAM8.DEC1.A_buf\[0\] SLICE\[0\].RAM8.DEC1.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[4\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_34_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[3\] BYTE\[2\].FLOATBUF0\[19\].Z Do0_REG.CLKBUF\[2\]
+ Do0[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_7_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_22_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_14_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_12_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_14_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_34_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_1_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_1_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[2\].W.SEL0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_27_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDEC1.AND3 A1BUF\[4\].X A1BUF\[3\].X DEC1.EN SLICE\[3\].RAM8.DEC1.EN VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_4_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_331 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_320 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_364 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_353 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_342 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[11\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[11\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_397 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_386 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_375 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND5 SLICE\[2\].RAM8.DEC0.A_buf_N\[1\] SLICE\[2\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[5\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_5_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_800 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_13_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X SLICE\[2\].RAM8.DEC0.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_32_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_25_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_1_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[18\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[18\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_27_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[0\].FLOATBUF0\[3\].__cell__ BYTE\[0\].FLOATBUF0\[3\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[3\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_18_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_11_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_26_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_11_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_24_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_7_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_652 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_641 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_630 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_696 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_685 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_674 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_663 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A SLICE\[2\].RAM8.WEBUF\[0\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_15_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.Root_CLKBUF CLKBUF.X Do0_REG.CLK_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_2_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_22_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_22_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.AND2 zero_ SLICE\[3\].RAM8.DEC1.A_buf_N\[0\] SLICE\[3\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[2\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_12_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_471 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_460 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_493 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A SLICE\[1\].RAM8.WEBUF\[2\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_17_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_17_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_21_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[7\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BYTE\[1\].FLOATBUF1\[12\].Z Do1_REG.CLKBUF\[1\]
+ Do1[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_14_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[1\].W.SEL0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_32_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[7\] BYTE\[3\].FLOATBUF0\[31\].Z Do0_REG.CLKBUF\[3\]
+ Do0[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_0_513 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_502 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC1.INV2 SLICE\[0\].RAM8.DEC1.A_buf\[1\] SLICE\[0\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_13_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_14_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_12_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_30_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_30_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_34_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_20_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_321 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_310 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_365 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_354 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_343 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_332 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_398 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_387 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_376 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[15\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[15\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XA0BUF\[1\].__cell__ A0[1] A0BUF\[1\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_3_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.DEC0.AND6 SLICE\[2\].RAM8.DEC0.A_buf_N\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[6\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_5_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_33_801 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_29_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_13_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_32_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_25_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_1_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_620 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_653 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_642 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_631 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_686 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_675 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_664 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_697 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_2_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_22_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF1\[21\].__cell__ BYTE\[2\].FLOATBUF1\[21\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[21\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.AND3 zero_ SLICE\[3\].RAM8.DEC1.A_buf\[1\] SLICE\[3\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[3\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\].X SLICE\[1\].RAM8.DEC1.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_12_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_20_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_2_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_28_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_17_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[3\].RAM8.WORD\[0\].W.SEL0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_33_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_33_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[4\] BYTE\[0\].FLOATBUF0\[4\].Z Do0_REG.CLKBUF\[0\]
+ Do0[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_4_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_0_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_25_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_16_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_28_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_16_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_32_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_0_514 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_503 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_18_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_4_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC1.INV3 SLICE\[0\].RAM8.DEC1.A_buf\[1\] SLICE\[0\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_7_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_22_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_30_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_1_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XTIE1\[1\].__cell__ BYTE\[1\].FLOATBUF1\[10\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xfill_27_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_20_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_29_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_322 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_311 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_300 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_355 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_344 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_333 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_399 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_388 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_377 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_366 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.AND7 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[2\].RAM8.DEC0.A_buf\[2\] SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.WORD\[7\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND0 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf_N SLICE\[0\].RAM8.WORD\[0\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xfill_13_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_25_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BYTE\[3\].FLOATBUF1\[25\].Z Do1_REG.CLKBUF\[3\]
+ Do1[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDIBUF\[3\].__cell__ Di0[3] DIBUF\[3\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_15_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF1\[3\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[3\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_8_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_610 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_643 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_632 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_621 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_687 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_676 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_665 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_654 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_698 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_30_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_26_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_9_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_2_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.AND4 SLICE\[3\].RAM8.DEC1.A_buf_N\[0\] SLICE\[3\].RAM8.DEC1.A_buf_N\[1\]
+ SLICE\[3\].RAM8.DEC1.A_buf\[2\] SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[4\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_12_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_462 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_495 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_484 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF1\[13\].__cell__ BYTE\[1\].FLOATBUF1\[13\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[13\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_20_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_28_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_33_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_21_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_4_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_0_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[7\].W.SEL0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_21_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_14_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_32_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_30_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_504 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_515 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC1.INV4 SLICE\[0\].RAM8.DEC1.EN_buf SLICE\[0\].RAM8.DEC1.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_34_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_22_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFBUFENBUF1\[1\].__cell__ EN1 BYTE\[1\].FLOATBUF1\[10\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_1_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_20_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_29_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_312 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_301 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_356 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_345 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_334 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_323 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_389 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_378 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_367 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[1\] BYTE\[2\].FLOATBUF0\[17\].Z Do0_REG.CLKBUF\[2\]
+ Do0[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_17_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND1 zero_ SLICE\[0\].RAM8.DEC0.A_buf_N\[1\] SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[1\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_25_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_18_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_15_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF1\[7\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[7\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_1_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_24_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_611 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_600 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_644 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_633 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_622 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_677 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_666 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_655 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X SLICE\[2\].RAM8.DEC0.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_699 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_688 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_30_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_23_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_26_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_30_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[31\].__cell__ BYTE\[3\].FLOATBUF0\[31\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[31\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF0\[2\].__cell__ BYTE\[0\].FLOATBUF0\[2\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[2\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.DEC1.AND5 SLICE\[3\].RAM8.DEC1.A_buf_N\[1\] SLICE\[3\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC1.A_buf\[2\] SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[5\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_12_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_485 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_2_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[6\].W.SEL0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_21_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_28_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_19_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_19_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[2\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[2\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_21_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_4_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_10_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_33_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[9\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[9\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_11_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_11_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_21_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_16_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_31_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[3\].FLOATBUF1\[26\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[26\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_505 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_516 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A SLICE\[1\].RAM8.WEBUF\[1\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_34_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_7_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_21_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BYTE\[1\].FLOATBUF1\[10\].Z Do1_REG.CLKBUF\[1\]
+ Do1[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_12_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_6_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.INV1 SLICE\[2\].RAM8.DEC0.A_buf\[0\] SLICE\[2\].RAM8.DEC0.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_1_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.CLKBUF.__cell__ CLKBUF.X SLICE\[3\].RAM8.CLKBUF.X VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_20_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_20_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_20_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[5\] BYTE\[3\].FLOATBUF0\[29\].Z Do0_REG.CLKBUF\[3\]
+ Do0[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_29_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_313 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_302 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_346 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_335 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_324 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_379 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_368 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_357 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\].X SLICE\[3\].RAM8.DEC1.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_17_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A SLICE\[0\].RAM8.WEBUF\[3\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_33_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_3_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_5_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_10_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_29_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND2 zero_ SLICE\[0\].RAM8.DEC0.A_buf_N\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[2\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_32_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_25_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_15_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_601 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_17_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_634 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_623 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_612 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_678 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_667 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_656 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_645 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_689 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_30_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[5\].W.SEL0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_23_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XA0BUF\[0\].__cell__ A0[0] A0BUF\[0\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_14_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_30_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC1.AND6 SLICE\[3\].RAM8.DEC1.A_buf_N\[0\] SLICE\[3\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC1.A_buf\[2\] SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[6\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_12_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[23\].__cell__ BYTE\[2\].FLOATBUF0\[23\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[23\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_464 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtap_21_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[3\].FLOATBUF1\[29\].__cell__ BYTE\[3\].FLOATBUF1\[29\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[29\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XBYTE\[1\].FLOATBUF0\[12\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[12\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_4_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[0\].FLOATBUF0\[6\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[6\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBYTE\[2\].FLOATBUF1\[23\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[23\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_23_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_21_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[19\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[19\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[20\].__cell__ BYTE\[2\].FLOATBUF1\[20\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[20\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_32_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[2\] BYTE\[0\].FLOATBUF0\[2\].Z Do0_REG.CLKBUF\[0\]
+ Do0[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_22_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_30_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_517 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_506 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_21_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BYTE\[2\].FLOATBUF1\[22\].Z Do1_REG.CLKBUF\[2\]
+ Do1[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_22_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.INV2 SLICE\[2\].RAM8.DEC0.A_buf\[1\] SLICE\[2\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_1_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XCLKBUF.__cell__ CLK CLKBUF.X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_1_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_20_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_4_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_29_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_303 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_347 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_336 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_325 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_314 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_369 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_358 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND3 zero_ SLICE\[0\].RAM8.DEC0.A_buf\[1\] SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[3\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_32_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[4\].W.SEL0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_25_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDIBUF\[29\].__cell__ Di0[29] DIBUF\[29\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_27_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.CLKBUF.__cell__ CLKBUF.X SLICE\[1\].RAM8.CLKBUF.X VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_28_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_28_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_18_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.ABUF\[2\] A1BUF\[2\].X SLICE\[0\].RAM8.DEC1.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_8_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTIE1\[0\].__cell__ BYTE\[0\].FLOATBUF1\[0\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_602 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_635 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_624 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_613 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_7_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_668 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_657 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_646 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_679 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_30_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_26_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[2\].__cell__ Di0[2] DIBUF\[2\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_14_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC1.AND7 SLICE\[3\].RAM8.DEC1.A_buf\[0\] SLICE\[3\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC1.A_buf\[2\] SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.WORD\[7\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_12_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_476 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_465 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_20_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.DEC1.AND0 SLICE\[1\].RAM8.DEC1.A_buf\[0\] SLICE\[1\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC1.A_buf\[2\] SLICE\[1\].RAM8.DEC1.EN_buf_N SLICE\[1\].RAM8.WORD\[0\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xfill_2_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtap_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[1\].FLOATBUF0\[15\].__cell__ BYTE\[1\].FLOATBUF0\[15\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[15\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_7_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_11_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_10_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_0_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_24_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XA1BUF\[4\].__cell__ A1[4] A1BUF\[4\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_8_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[6\] BYTE\[1\].FLOATBUF0\[14\].Z Do0_REG.CLKBUF\[1\]
+ Do0[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[12\].__cell__ BYTE\[1\].FLOATBUF1\[12\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[12\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_18_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_518 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_0_507 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDEC1.INV1 A1BUF\[3\].X DEC1.A_N\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_7_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_21_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[1\].FLOATBUF0\[9\].__cell__ BYTE\[1\].FLOATBUF0\[9\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[9\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_12_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[3\].W.SEL0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_6_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.INV3 SLICE\[2\].RAM8.DEC0.A_buf\[1\] SLICE\[2\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[19\].__cell__ Di0[19] DIBUF\[19\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xtap_1_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_29_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_304 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_337 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_326 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_315 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_359 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_348 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_5_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.AND4 SLICE\[0\].RAM8.DEC0.A_buf_N\[0\] SLICE\[0\].RAM8.DEC0.A_buf_N\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[4\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_25_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_18_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFBUFENBUF1\[0\].__cell__ EN1 BYTE\[0\].FLOATBUF1\[0\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_26_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_625 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_614 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_603 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_669 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_658 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_647 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_636 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_30_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_31_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_30_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_2_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_12_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_12_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_499 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_20_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.AND1 zero_ SLICE\[1\].RAM8.DEC1.A_buf_N\[1\] SLICE\[1\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[1\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BYTE\[0\].FLOATBUF1\[7\].Z Do1_REG.CLKBUF\[0\]
+ Do1[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_0_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[3\].FLOATBUF0\[30\].__cell__ BYTE\[3\].FLOATBUF0\[30\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[30\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[2\].W.SEL0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_8_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[1\].__cell__ BYTE\[0\].FLOATBUF0\[1\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[1\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_19_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_30_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_9_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_519 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_508 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_18_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDEC1.INV2 A1BUF\[4\].X DEC1.A_N\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_12_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.INV4 SLICE\[2\].RAM8.DEC0.EN_buf SLICE\[2\].RAM8.DEC0.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_20_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_29_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_338 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_327 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_316 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_305 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_349 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X SLICE\[1\].RAM8.DEC0.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_3_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BYTE\[1\].FLOATBUF1\[8\].Z Do1_REG.CLKBUF\[1\]
+ Do1[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_29_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND5 SLICE\[0\].RAM8.DEC0.A_buf_N\[1\] SLICE\[0\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[5\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A SLICE\[1\].RAM8.WEBUF\[0\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_18_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_15_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[3\] BYTE\[3\].FLOATBUF0\[27\].Z Do0_REG.CLKBUF\[3\]
+ Do0[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_28_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.Root_CLKBUF CLKBUF.X Do1_REG.CLK_buf VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_26_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_626 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_615 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_604 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_659 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_648 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_637 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_30_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_16_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WEBUF\[2\].__cell__ SLICE\[0\].RAM8.WEBUF\[2\].A SLICE\[0\].RAM8.WEBUF\[2\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_9_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.DEC1.INV1 SLICE\[3\].RAM8.DEC1.A_buf\[0\] SLICE\[3\].RAM8.DEC1.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_30_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_12_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_12_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.AND2 zero_ SLICE\[1\].RAM8.DEC1.A_buf_N\[0\] SLICE\[1\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[2\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_21_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[1\].W.SEL0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_11_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_0_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_25_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_16_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF0\[22\].__cell__ BYTE\[2\].FLOATBUF0\[22\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[22\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[3\].FLOATBUF1\[28\].__cell__ BYTE\[3\].FLOATBUF1\[28\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[28\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_15_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_509 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_18_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDEC1.INV3 DEC1.EN DEC1.EN_N VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_12_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_1_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_31_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[0\] BYTE\[0\].FLOATBUF0\[0\].Z Do0_REG.CLKBUF\[0\]
+ Do0[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_20_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_29_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_328 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_317 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_306 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_339 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_17_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BYTE\[2\].FLOATBUF1\[20\].Z Do1_REG.CLKBUF\[2\]
+ Do1[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_3_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_29_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC0.AND0 A0BUF\[3\].X A0BUF\[4\].X DEC0.EN_N SLICE\[0\].RAM8.DEC0.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xfill_29_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND6 SLICE\[0\].RAM8.DEC0.A_buf_N\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[6\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_15_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[7\].W.SEL1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_31_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[2\].FLOATBUF0\[20\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[20\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_28_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[3\].FLOATBUF1\[31\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[31\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_17_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_616 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_605 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_7_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_7_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_649 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_638 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_627 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_30_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[3\].FLOATBUF0\[27\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[27\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_16_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_26_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.DEC1.INV2 SLICE\[3\].RAM8.DEC1.A_buf\[1\] SLICE\[3\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_9_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[2\].RAM8.WORD\[0\].W.SEL0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_14_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC1.ABUF\[0\] A1BUF\[0\].X SLICE\[0\].RAM8.DEC1.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDIBUF\[28\].__cell__ Di0[28] DIBUF\[28\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_14_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_435 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_424 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_413 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_402 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_468 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_457 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_446 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_479 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.AND3 zero_ SLICE\[1\].RAM8.DEC1.A_buf\[1\] SLICE\[1\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[3\].W.SEL1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xtap_21_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_14_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_7_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_28_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_4_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_4_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_10_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_276 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_265 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_254 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_298 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_287 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_11_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[1\].__cell__ Di0[1] DIBUF\[1\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_5_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XTIE0\[3\].__cell__ BYTE\[3\].FLOATBUF0\[24\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_8_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_8_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_26_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[10\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[10\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[14\].__cell__ BYTE\[1\].FLOATBUF0\[14\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[14\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_15_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_9_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_18_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_12_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[2\].FLOATBUF1\[17\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[17\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_1_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[4\] BYTE\[1\].FLOATBUF0\[12\].Z Do0_REG.CLKBUF\[1\]
+ Do0[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_24_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[6\].W.SEL1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_20_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_29_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_329 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_318 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_307 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XA1BUF\[3\].__cell__ A1[3] A1BUF\[3\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_17_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_3_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[11\].__cell__ BYTE\[1\].FLOATBUF1\[11\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[11\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC0.AND1 DEC0.A_N\[1\] A0BUF\[3\].X DEC0.EN SLICE\[1\].RAM8.DEC0.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
Xfill_29_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.AND7 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[0\].RAM8.DEC0.A_buf\[2\] SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.WORD\[7\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_15_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_2_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF0\[8\].__cell__ BYTE\[1\].FLOATBUF0\[8\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[8\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[18\].__cell__ Di0[18] DIBUF\[18\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_8_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_17_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_7_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_617 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_606 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_7_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_639 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_628 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_23_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.DEC1.INV3 SLICE\[3\].RAM8.DEC1.A_buf\[1\] SLICE\[3\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_9_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_14_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_30_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_22_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_490 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_425 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_414 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_403 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[7\].W.SEL0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_12_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_458 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_447 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_436 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_469 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC1.AND4 SLICE\[1\].RAM8.DEC1.A_buf_N\[0\] SLICE\[1\].RAM8.DEC1.A_buf_N\[1\]
+ SLICE\[1\].RAM8.DEC1.A_buf\[2\] SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[4\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_21_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_7_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_28_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[3\].RAM8.DEC0.AND0 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf_N SLICE\[3\].RAM8.WORD\[0\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xtap_4_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_10_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_23_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_23_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_277 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_266 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_255 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_299 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_288 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_11_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_5_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFBUFENBUF0\[3\].__cell__ EN0 BYTE\[3\].FLOATBUF0\[24\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_244 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_8_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[5\].W.SEL1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[14\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[14\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_15_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF1\[7\].__cell__ BYTE\[0\].FLOATBUF1\[7\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[7\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_30_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BYTE\[0\].FLOATBUF1\[5\].Z Do1_REG.CLKBUF\[0\]
+ Do1[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_18_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_6_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_17_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_20_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_29_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_319 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_308 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[0\].__cell__ BYTE\[0\].FLOATBUF0\[0\].TE_BN BYTE\[0\].FLOATBUF0\[0\].A
+ BYTE\[0\].FLOATBUF0\[0\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_3_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC0.AND2 DEC0.A_N\[0\] A0BUF\[4\].X DEC0.EN SLICE\[2\].RAM8.DEC0.EN VDD VDD VSS
+ VSS gf180mcu_fd_sc_mcu7t5v0__and3_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_15_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_2_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_8_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X SLICE\[1\].RAM8.DEC0.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_607 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[6\].W.SEL0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_7_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_629 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_618 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_17_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.DEC1.INV4 SLICE\[3\].RAM8.DEC1.EN_buf SLICE\[3\].RAM8.DEC1.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_9_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_14_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[3\].Do_FF\[1\] BYTE\[3\].FLOATBUF0\[25\].Z Do0_REG.CLKBUF\[3\]
+ Do0[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_31_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_491 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_480 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_426 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_415 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_404 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_12_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_459 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_448 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_437 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_20_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.AND5 SLICE\[1\].RAM8.DEC1.A_buf_N\[1\] SLICE\[1\].RAM8.DEC1.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC1.A_buf\[2\] SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[5\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_21_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_7_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_25_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_11_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[4\].W.SEL1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_28_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC0.AND1 zero_ SLICE\[3\].RAM8.DEC0.A_buf_N\[1\] SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[1\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[0\].RAM8.WEBUF\[1\].__cell__ SLICE\[0\].RAM8.WEBUF\[1\].A SLICE\[0\].RAM8.WEBUF\[1\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_15_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_10_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_267 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_256 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_289 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_278 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_24_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_245 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_790 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_9_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_30_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_18_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_18_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_22_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_6_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[0\].FLOATBUF1\[2\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[2\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.INV1 SLICE\[0\].RAM8.DEC0.A_buf\[0\] SLICE\[0\].RAM8.DEC0.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_24_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_17_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\].X SLICE\[2\].RAM8.DEC1.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_0_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_20_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_9_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_309 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[9\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[9\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[21\].__cell__ BYTE\[2\].FLOATBUF0\[21\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[21\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.Do_CLKBUF\[2\] Do1_REG.CLK_buf Do1_REG.CLKBUF\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_33_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_10_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[27\].__cell__ BYTE\[3\].FLOATBUF1\[27\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[27\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[3\].DIODE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_5_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDEC0.AND3 A0BUF\[4\].X A0BUF\[3\].X DEC0.EN SLICE\[3\].RAM8.DEC0.EN VDD VDD VSS VSS
+ gf180mcu_fd_sc_mcu7t5v0__and3_2
XSLICE\[1\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[5\].W.SEL0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_23_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_15_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BYTE\[2\].FLOATBUF1\[18\].Z Do1_REG.CLKBUF\[2\]
+ Do1[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_608 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_17_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_619 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_26_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_9_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[3\].W.SEL1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_22_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_492 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_481 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_470 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_12_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_416 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_405 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_12_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_449 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_438 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_427 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC1.ENBUF SLICE\[2\].RAM8.DEC1.EN SLICE\[2\].RAM8.DEC1.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_13_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.DEC1.AND6 SLICE\[1\].RAM8.DEC1.A_buf_N\[0\] SLICE\[1\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC1.A_buf\[2\] SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[6\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_14_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_27_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC0.AND2 zero_ SLICE\[3\].RAM8.DEC0.A_buf_N\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[2\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_15_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_3_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_3_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_23_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_18_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_268 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_257 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_279 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDIBUF\[27\].__cell__ Di0[27] DIBUF\[27\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xtap_12_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_246 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_24_235 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_780 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_791 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_9_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_30_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtap_18_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_18_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[4\].W.SEL0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBYTE\[0\].FLOATBUF1\[6\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[6\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.INV2 SLICE\[0\].RAM8.DEC0.A_buf\[1\] SLICE\[0\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[2\].DIODE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_24_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_0_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_20_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[0\].__cell__ Di0[0] DIBUF\[0\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_9_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_9_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XTIE0\[2\].__cell__ BYTE\[2\].FLOATBUF0\[16\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_17_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_33_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_10_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XBYTE\[1\].FLOATBUF0\[13\].__cell__ BYTE\[1\].FLOATBUF0\[13\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[13\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF1\[19\].__cell__ BYTE\[2\].FLOATBUF1\[19\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[19\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[2\] BYTE\[1\].FLOATBUF0\[10\].Z Do0_REG.CLKBUF\[1\]
+ Do0[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_2_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_15_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_22_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_2_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_58 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[2\].W.SEL1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[6\] BYTE\[3\].FLOATBUF1\[30\].Z Do1_REG.CLKBUF\[3\]
+ Do1[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_28_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_26_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_26_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_18_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_609 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XA1BUF\[2\].__cell__ A1[2] A1BUF\[2\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_25_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[1\].FLOATBUF1\[10\].__cell__ BYTE\[1\].FLOATBUF1\[10\].TE_BN BYTE\[1\].FLOATBUF1\[10\].A
+ BYTE\[1\].FLOATBUF1\[10\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[1\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[1\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_14_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_22_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XBYTE\[1\].FLOATBUF0\[8\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[8\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_20_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_482 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_471 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_460 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_90 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_493 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_12_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_417 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_406 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_439 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_428 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_13_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.AND7 SLICE\[1\].RAM8.DEC1.A_buf\[0\] SLICE\[1\].RAM8.DEC1.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC1.A_buf\[2\] SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.WORD\[7\].W.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_13_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_21_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[17\].__cell__ Di0[17] DIBUF\[17\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xtap_14_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[3\].FLOATBUF1\[25\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[25\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_7_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_8_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_33_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_233 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_27_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.AND3 zero_ SLICE\[3\].RAM8.DEC0.A_buf\[1\] SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[3\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_15_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_290 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_23_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_23_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_258 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_269 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_11_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_12_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_5_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[3\].W.SEL0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_13_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_247 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_236 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_781 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_770 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_792 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_8_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.ENBUF SLICE\[2\].RAM8.DEC0.EN SLICE\[2\].RAM8.DEC0.EN_buf VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_26_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_19_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X SLICE\[3\].RAM8.DEC0.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_18_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_18_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_34_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_34_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_22_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_21_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_6_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.INV3 SLICE\[0\].RAM8.DEC0.A_buf\[1\] SLICE\[0\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[0\].W.CLKBUF SLICE\[1\].RAM8.CLKBUF.X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_24_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_17_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF1\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_20_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF0\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFBUFENBUF0\[2\].__cell__ EN0 BYTE\[2\].FLOATBUF0\[16\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_9_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_9_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_29_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[3\] BYTE\[0\].FLOATBUF1\[3\].Z Do1_REG.CLKBUF\[0\]
+ Do1[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[3\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[1\].W.SEL1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_19_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_5_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF1\[6\].__cell__ BYTE\[0\].FLOATBUF1\[6\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[6\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[6\] BYTE\[2\].FLOATBUF0\[22\].Z Do0_REG.CLKBUF\[2\]
+ Do0[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_29_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF1\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_15_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_22_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_15_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_31_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_18_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_32_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_6_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[11\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[11\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_31_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF0\[5\].TE_BINV BYTE\[0\].FLOATBUF0\[0\].TE_B BYTE\[0\].FLOATBUF0\[5\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_28_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[2\].FLOATBUF1\[22\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[22\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_16_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_32_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_450 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_483 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_472 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_461 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_494 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_91 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_407 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_429 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_418 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBYTE\[2\].FLOATBUF0\[18\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[18\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_14_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_7_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[2\].W.SEL0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_25_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[29\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[29\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_25_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_26_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_27_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_234 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_15_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.AND4 SLICE\[3\].RAM8.DEC0.A_buf_N\[0\] SLICE\[3\].RAM8.DEC0.A_buf_N\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[4\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_15_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_10_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_291 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_280 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_23_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_2_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_18_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_259 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_11_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_5_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_13_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_248 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_24_237 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_771 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_760 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1INV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_793 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_782 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_30_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.SEL1BUF SLICE\[3\].RAM8.WORD\[0\].W.SEL1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_18_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_34_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_34_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[3\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_5_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WEBUF\[0\].__cell__ SLICE\[0\].RAM8.WEBUF\[0\].A SLICE\[0\].RAM8.WEBUF\[0\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_10_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_12_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_33_590 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_24_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.DEC0.INV4 SLICE\[0\].RAM8.DEC0.EN_buf SLICE\[0\].RAM8.DEC0.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[7\] BYTE\[1\].FLOATBUF1\[15\].Z Do1_REG.CLKBUF\[1\]
+ Do1[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_17_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[2\] BYTE\[1\].FLOATBUF1\[10\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.ABUF\[2\] A0BUF\[2\].X SLICE\[0\].RAM8.DEC0.A_buf\[2\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_9_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XEN1BUF.__cell__ EN1 DEC1.EN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_5_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_19_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF0\[29\].__cell__ BYTE\[3\].FLOATBUF0\[29\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[29\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_23_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_2_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_31_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_0_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_2_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_49 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.Do_CLKBUF\[0\] Do1_REG.CLK_buf Do1_REG.CLKBUF\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_21_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.CGAND SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[0\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_17_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_17_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_6_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF0\[20\].__cell__ BYTE\[2\].FLOATBUF0\[20\].TE_BN BYTE\[2\].FLOATBUF0\[16\].A
+ BYTE\[2\].FLOATBUF0\[20\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_6_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[1\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[1\].W.SEL0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XBYTE\[3\].FLOATBUF1\[26\].__cell__ BYTE\[3\].FLOATBUF1\[26\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[26\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[15\].TE_BINV BYTE\[1\].FLOATBUF0\[10\].TE_B BYTE\[1\].FLOATBUF0\[15\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_14_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.INV1 SLICE\[1\].RAM8.DEC1.A_buf\[0\] SLICE\[1\].RAM8.DEC1.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].Do_FF\[0\] BYTE\[2\].FLOATBUF1\[16\].Z Do1_REG.CLKBUF\[2\]
+ Do1[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_22_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_440 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_473 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_462 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_451 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_495 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_484 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_92 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_408 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_419 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_7_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_8_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtap_26_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_15_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.AND5 SLICE\[3\].RAM8.DEC0.A_buf_N\[1\] SLICE\[3\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[5\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_15_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_31_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_0_292 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_281 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_270 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_11_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_12_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_13_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_249 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_24_238 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_772 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_761 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_750 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_794 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_783 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_26_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_15_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_15_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XEN0BUF.__cell__ EN0 DEC0.EN VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_34_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[7\] BYTE\[0\].FLOATBUF0\[7\].Z Do0_REG.CLKBUF\[0\]
+ Do0[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_22_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_21_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_10_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_3_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_580 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_33_591 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_12_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[7\].W.SEL1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[26\].__cell__ Di0[26] DIBUF\[26\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_0_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_29_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_17_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_3_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_19_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_1_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.SEL0BUF SLICE\[1\].RAM8.WORD\[0\].W.SEL0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_28_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTIE0\[1\].__cell__ BYTE\[1\].FLOATBUF0\[10\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].Do_FF\[0\] BYTE\[1\].FLOATBUF0\[8\].Z Do0_REG.CLKBUF\[1\]
+ Do0[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_6_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF0\[12\].__cell__ BYTE\[1\].FLOATBUF0\[12\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[12\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC1.INV2 SLICE\[1\].RAM8.DEC1.A_buf\[1\] SLICE\[1\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF1\[18\].__cell__ BYTE\[2\].FLOATBUF1\[18\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[18\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_28_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[4\] BYTE\[3\].FLOATBUF1\[28\].Z Do1_REG.CLKBUF\[3\]
+ Do1[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_32_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_22_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_4_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_20_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_441 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_430 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_474 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_463 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_452 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_71 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_60 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_496 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_485 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_93 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_82 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[3\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_33_409 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_25_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_33_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_19_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XA1BUF\[1\].__cell__ A1[1] A1BUF\[1\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.AND6 SLICE\[3\].RAM8.DEC0.A_buf_N\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[6\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_15_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_282 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_271 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_260 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_293 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_33_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[2\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_12_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_5_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_239 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_762 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_751 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_740 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_33_795 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_784 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_773 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_31_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[6\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[6\].W.SEL1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDIBUF\[16\].__cell__ Di0[16] DIBUF\[16\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_9_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_5_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_5_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[1\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_10_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_3_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_570 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_592 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_581 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_12_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_5_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[1\].DIODE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_17_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_10_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_3_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_19_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_19_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_1_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_2_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_15_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.Do_CLKBUF\[2\] Do0_REG.CLK_buf Do0_REG.CLKBUF\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_28_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_28_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_2_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo1_REG.OUTREG_BYTE\[0\].Do_FF\[1\] BYTE\[0\].FLOATBUF1\[1\].Z Do1_REG.CLKBUF\[0\]
+ Do1[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_28_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_26_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF0\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[7\].W.SEL0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_18_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFBUFENBUF0\[1\].__cell__ EN0 BYTE\[1\].FLOATBUF0\[10\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_18_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[4\] BYTE\[2\].FLOATBUF0\[20\].Z Do0_REG.CLKBUF\[2\]
+ Do0[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_17_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_7_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_6_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[0\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_13_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_16_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC1.INV3 SLICE\[1\].RAM8.DEC1.A_buf\[1\] SLICE\[1\].RAM8.DEC1.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XBYTE\[0\].FLOATBUF1\[5\].__cell__ BYTE\[0\].FLOATBUF1\[5\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[5\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_16_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_32_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_431 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_420 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_464 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_453 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_442 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_50 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_497 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_486 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_475 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_94 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_4_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_25_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[5\].W.SEL1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_33_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_1_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtap_26_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.AND7 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[3\].RAM8.DEC0.A_buf\[2\] SLICE\[3\].RAM8.DEC0.EN_buf SLICE\[3\].RAM8.WORD\[7\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_15_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_10_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.DEC0.AND0 SLICE\[1\].RAM8.DEC0.A_buf\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.A_buf\[2\] SLICE\[1\].RAM8.DEC0.EN_buf_N SLICE\[1\].RAM8.WORD\[0\].W.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xfill_10_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].genblk1.STORAGE DIBUF\[5\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_283 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_272 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_261 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_250 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_294 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_226 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_18_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_12_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_5_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_13_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_24_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_763 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_752 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_741 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_730 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_796 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_785 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_774 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_32_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_31_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_15_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_23_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_5_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].genblk1.STORAGE DIBUF\[22\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_5_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_24_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_3_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDo0_REG.OUTREG_BYTE\[0\].DIODE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_571 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_560 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_593 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_582 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_6_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDEC0.INV1 A0BUF\[3\].X DEC0.A_N\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[2\].DIODE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_9_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[30\].TE_BINV BYTE\[3\].FLOATBUF1\[24\].TE_B BYTE\[3\].FLOATBUF1\[30\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_5_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[2\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.CLKBUF SLICE\[0\].RAM8.CLKBUF.X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_10_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_3_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_19_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[6\].W.SEL0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XBYTE\[3\].FLOATBUF0\[26\].TE_BINV BYTE\[3\].FLOATBUF0\[24\].TE_B BYTE\[3\].FLOATBUF0\[26\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_29_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[6\].genblk1.STORAGE DIBUF\[30\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_29_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.CGAND SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[3\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF0\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[5\].genblk1.STORAGE DIBUF\[13\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_390 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XDo1_REG.OUTREG_BYTE\[1\].Do_FF\[5\] BYTE\[1\].FLOATBUF1\[13\].Z Do1_REG.CLKBUF\[1\]
+ Do1[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_15_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_28_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.DEC0.ABUF\[0\] A0BUF\[0\].X SLICE\[0\].RAM8.DEC0.A_buf\[0\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_2_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_2_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_21_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[5\] BYTE\[2\].FLOATBUF1\[21\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF0\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_18_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[2\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_25_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_6_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].genblk1.STORAGE DIBUF\[4\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_16_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[0\].genblk1.STORAGE DIBUF\[16\].X SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_16_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC1.INV4 SLICE\[1\].RAM8.DEC1.EN_buf SLICE\[1\].RAM8.DEC1.EN_buf_N
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XBYTE\[3\].FLOATBUF0\[28\].__cell__ BYTE\[3\].FLOATBUF0\[28\].TE_BN BYTE\[3\].FLOATBUF0\[24\].A
+ BYTE\[3\].FLOATBUF0\[28\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[4\].W.SEL1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_28_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_204 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_215 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_20_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_432 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_421 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_410 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_465 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_454 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_443 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_51 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_498 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_487 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_476 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_73 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_102 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_124 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[1\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_13_157 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_168 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_179 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_21_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_8_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_33_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_12_190 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_27_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[5\].genblk1.STORAGE DIBUF\[21\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_27_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_27_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_31_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[2\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_10_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.DEC0.AND1 zero_ SLICE\[1\].RAM8.DEC0.A_buf_N\[1\] SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[1\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
Xfill_10_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[3\].FLOATBUF1\[25\].__cell__ BYTE\[3\].FLOATBUF1\[25\].TE_BN BYTE\[3\].FLOATBUF1\[24\].A
+ BYTE\[3\].FLOATBUF1\[25\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_240 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_273 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_262 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_251 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_295 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_284 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_227 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_18_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[2\].FLOATBUF1\[16\].TE_BINV BYTE\[2\].FLOATBUF1\[16\].TE_B BYTE\[2\].FLOATBUF1\[16\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_5_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_720 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_753 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_742 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_731 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_786 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_775 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_764 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_797 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtap_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_219 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[5\].genblk1.STORAGE DIBUF\[29\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[5\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_23_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[4\].genblk1.STORAGE DIBUF\[12\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[0\].genblk1.STORAGE DIBUF\[24\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtap_5_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_5_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[1\].DIODE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[5\].W.SEL0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_10_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[3\].W.CLKBUF SLICE\[3\].RAM8.CLKBUF.X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xtap_3_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_24_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.DEC1.ABUF\[1\] A1BUF\[1\].X SLICE\[1\].RAM8.DEC1.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_561 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_550 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_594 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_583 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_572 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_222 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XBYTE\[2\].FLOATBUF0\[23\].TE_BINV BYTE\[2\].FLOATBUF0\[16\].TE_B BYTE\[2\].FLOATBUF0\[23\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDEC0.INV2 A0BUF\[4\].X DEC0.A_N\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[2\].RAM8.WEBUF\[0\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_24_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_17_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_200 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_211 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_5_140 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_162 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_173 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_184 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_195 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[4\].genblk1.STORAGE DIBUF\[20\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo0_REG.OUTREG_BYTE\[0\].Do_FF\[5\] BYTE\[0\].FLOATBUF0\[5\].Z Do0_REG.CLKBUF\[0\]
+ Do0[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtap_10_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].genblk1.STORAGE DIBUF\[3\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_10_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_1_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_29_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[1\] BYTE\[2\].FLOATBUF1\[17\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF0 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF0\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_23_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_380 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_391 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_132 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_110 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_165 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_154 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.genblk1.CG SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.CLK_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.WE0_WIRE
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_2_198 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_187 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_176 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xfill_28_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[3\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[3\].W.SEL1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_2_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_19_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_21_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[6\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[6\] BYTE\[0\].FLOATBUF1\[6\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDIBUF\[25\].__cell__ Di0[25] DIBUF\[25\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF0\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_202 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_213 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_224 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_28_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_16_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_32_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_22_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_205 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_216 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfill_30_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_422 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_411 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_400 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_455 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_444 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_433 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_52 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_499 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_488 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_477 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_466 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_96 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.DEC0.INV1 SLICE\[3\].RAM8.DEC0.A_buf\[0\] SLICE\[3\].RAM8.DEC0.A_buf_N\[0\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF0\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_13_158 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_169 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF0\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_21_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[4\].genblk1.STORAGE DIBUF\[28\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[4\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[3\].genblk1.STORAGE DIBUF\[11\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDIBUF\[9\].__cell__ Di0[9] DIBUF\[9\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfill_9_1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XBYTE\[1\].FLOATBUF1\[13\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[13\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_33_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_1_208 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_12_180 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_191 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTIE0\[0\].__cell__ BYTE\[0\].FLOATBUF0\[0\].A VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xtap_26_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XDo1_REG.OUTREG_BYTE\[3\].Do_FF\[2\] BYTE\[3\].FLOATBUF1\[26\].Z Do1_REG.CLKBUF\[3\]
+ Do1[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfill_27_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_228 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF1\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF0\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF0\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC0.AND2 zero_ SLICE\[1\].RAM8.DEC0.A_buf_N\[0\] SLICE\[1\].RAM8.DEC0.A_buf\[1\]
+ SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[2\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XBYTE\[1\].FLOATBUF0\[11\].__cell__ BYTE\[1\].FLOATBUF0\[11\].TE_BN BYTE\[1\].FLOATBUF0\[10\].A
+ BYTE\[1\].FLOATBUF0\[11\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_230 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF1\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_274 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_263 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_252 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_241 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF0\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_296 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_285 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_3_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[2\].FLOATBUF1\[17\].__cell__ BYTE\[2\].FLOATBUF1\[17\].TE_BN BYTE\[2\].FLOATBUF1\[16\].A
+ BYTE\[2\].FLOATBUF1\[17\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_18_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_18_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF0\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_33_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[4\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[4\].W.SEL0 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XSLICE\[2\].RAM8.WORD\[6\].W.CLKBUF SLICE\[2\].RAM8.CLKBUF.X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[0\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF1\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF0 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF0\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_710 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_24_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_754 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_743 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_732 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_721 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_33_787 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_776 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_765 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_798 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo1_REG.OUTREG_BYTE\[0\].DIODE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF1\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[3\].genblk1.STORAGE DIBUF\[19\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_31_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF1\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_17_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[2\].genblk1.STORAGE DIBUF\[2\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.DIODE_CLK SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_26_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_209 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_105 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_116 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_127 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_149 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_23_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF1\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_14_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XA1BUF\[0\].__cell__ A1[0] A1BUF\[0\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_5_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_5_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_160 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_171 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_182 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_193 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[5\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF1\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0INV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_3_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_24_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.CGAND SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[2\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_33_562 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_551 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_540 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF1\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_6_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_595 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_584 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_573 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_223 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfill_12_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[2\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF0\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDEC0.INV3 DEC0.EN DEC0.EN_N VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_17_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_0_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[2\].genblk1.STORAGE DIBUF\[10\].X SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[2\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[2\].W.SEL1 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_9_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_201 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_212 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_5_152 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_163 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_174 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_5_185 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_5_196 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_10_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[3\].B.DIODE_CLK SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_19_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XDIBUF\[15\].__cell__ Di0[15] DIBUF\[15\].X VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_1_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_29_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.BIT\[6\].OBUF1 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF1\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[2\].OBUF1 SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[2\] BYTE\[0\].FLOATBUF1\[2\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[1\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF0\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_23_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_370 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_23_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_392 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_381 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.CGAND SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[1\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].OBUF0 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF0\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_2_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_111 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_100 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_166 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_155 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_199 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_188 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_2_177 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_28_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_28_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.CGAND SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[3\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtap_2_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_2_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF1\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[3\].genblk1.STORAGE DIBUF\[27\].X SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[3\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_19_120 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_153 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF0\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_21_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_19_197 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_186 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_175 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_19_164 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xtap_21_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_21_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.genblk1.CLKINV SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[5\].OBUF1 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[5\] BYTE\[3\].FLOATBUF1\[29\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[6\] BYTE\[1\].FLOATBUF0\[14\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.BIT\[7\].OBUF1 SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF1\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_18_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0INV SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[2\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_25_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_25_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_203 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_7_214 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.OUTREG_BYTE\[3\].DIODE\[1\] BYTE\[3\].FLOATBUF0\[25\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].genblk1.STORAGE DIBUF\[7\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_7_225 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_56 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_67 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_78 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_6_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[4\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_20_4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[0\] BYTE\[2\].FLOATBUF0\[16\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XDo0_REG.Do_CLKBUF\[0\] Do0_REG.CLK_buf Do0_REG.CLKBUF\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfill_16_112 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_145 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_16_189 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_178 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_167 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_16_156 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.BIT\[0\].genblk1.STORAGE DIBUF\[0\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[0\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1INV SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_28_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF1\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.CGAND SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WEBUF\[1\].X SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[1\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.DIODE_CLK SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xtap_16_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_16_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_22_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.genblk1.CG SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.CLK_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.WE0_WIRE
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[3\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_22_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_22_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_22_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[7\].genblk1.STORAGE DIBUF\[23\].X SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_4_206 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_4_217 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfill_30_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_30_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_20_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_423 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_412 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_401 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_456 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_445 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_434 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_489 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_478 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_467 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_86 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_75 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_29_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].genblk1.STORAGE DIBUF\[18\].X SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[0\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[0\] BYTE\[3\].FLOATBUF0\[24\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.DEC0.INV2 SLICE\[3\].RAM8.DEC0.A_buf\[1\] SLICE\[3\].RAM8.DEC0.A_buf_N\[1\]
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[1\].genblk1.STORAGE DIBUF\[1\].X SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XDo0_REG.OUTREG_BYTE\[2\].Do_FF\[2\] BYTE\[2\].FLOATBUF0\[18\].Z Do0_REG.CLKBUF\[2\]
+ Do0[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[2\] BYTE\[2\].FLOATBUF1\[18\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[3\] BYTE\[0\].FLOATBUF0\[3\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_13_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_126 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_13_159 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[3\].W.SEL0BUF SLICE\[0\].RAM8.WORD\[3\].W.SEL0 SLICE\[0\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_21_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_21_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[2\].B.Q_WIRE\[4\] BYTE\[2\].FLOATBUF1\[20\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[3\].W.BYTE\[0\].B.Q_WIRE\[5\] BYTE\[0\].FLOATBUF0\[5\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_9_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_11_0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_8_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_8_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[1\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XFBUFENBUF0\[0\].__cell__ EN0 BYTE\[0\].FLOATBUF0\[0\].TE_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_12_170 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_33_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_12_181 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_12_192 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_26_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[2\].W.BYTE\[2\].B.Q_WIRE\[7\] BYTE\[2\].FLOATBUF0\[23\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_1_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_19_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_27_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.CGAND SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL0
+ SLICE\[1\].RAM8.WEBUF\[0\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[0\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_27_229 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_27_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[1\].genblk1.STORAGE DIBUF\[17\].X SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_15_33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_66 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_55 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] BYTE\[3\].FLOATBUF1\[26\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[1\] BYTE\[0\].FLOATBUF1\[1\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_15_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_88 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_15_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[3\].OBUF0 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[3\] BYTE\[1\].FLOATBUF0\[11\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_31_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.genblk1.CLKINV SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[3\].B.CLK_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_10_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_10_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_31_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[4\].OBUF1 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[4\] BYTE\[3\].FLOATBUF1\[28\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.BIT\[5\].OBUF0 SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[3\].RAM8.WORD\[6\].W.BYTE\[1\].B.Q_WIRE\[5\] BYTE\[1\].FLOATBUF0\[13\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.DEC0.AND3 zero_ SLICE\[1\].RAM8.DEC0.A_buf\[1\] SLICE\[1\].RAM8.DEC0.A_buf\[0\]
+ SLICE\[1\].RAM8.DEC0.EN_buf SLICE\[1\].RAM8.WORD\[3\].W.SEL0 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and4_2
XSLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.CGAND SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL0
+ SLICE\[3\].RAM8.WEBUF\[2\].X SLICE\[3\].RAM8.WORD\[0\].W.BYTE\[2\].B.WE0_WIRE VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfill_0_231 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_220 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.genblk1.CG SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.CLK_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xfill_0_264 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_253 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_242 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[0\].FLOATBUF1\[4\].__cell__ BYTE\[0\].FLOATBUF1\[4\].TE_BN BYTE\[0\].FLOATBUF1\[0\].A
+ BYTE\[0\].FLOATBUF1\[4\].Z VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[2\].W.BYTE\[0\].B.Q_WIRE\[7\] BYTE\[0\].FLOATBUF1\[7\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_0_297 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_286 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_0_275 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_57 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.BIT\[7\].genblk1.STORAGE DIBUF\[31\].X SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[6\].W.BYTE\[3\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_2_9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_3_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_218 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_18_207 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[2\].B.Q_WIRE\[3\] BYTE\[2\].FLOATBUF1\[19\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[6\].genblk1.STORAGE DIBUF\[14\].X SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.GCLK
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.Q_WIRE\[4\] BYTE\[0\].FLOATBUF0\[4\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[2\].genblk1.STORAGE DIBUF\[26\].X SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[2\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.BIT\[7\].OBUF0 SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[5\].W.BYTE\[3\].B.Q_WIRE\[7\] BYTE\[3\].FLOATBUF0\[31\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[1\].genblk1.STORAGE DIBUF\[9\].X SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.GCLK
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[1\].RAM8.WORD\[2\].W.BYTE\[1\].B.DIODE_CLK SLICE\[1\].RAM8.WORD\[2\].W.BYTE\[0\].B.CLK
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XBYTE\[0\].FLOATBUF1\[1\].TE_BINV BYTE\[0\].FLOATBUF1\[0\].TE_B BYTE\[0\].FLOATBUF1\[1\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_13_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1INV SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL1
+ SLICE\[3\].RAM8.WORD\[7\].W.BYTE\[1\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[1\].OBUF1 SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[1\] BYTE\[1\].FLOATBUF1\[9\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[0\].W.BYTE\[2\].B.Q_WIRE\[6\] BYTE\[2\].FLOATBUF0\[22\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_13_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_13_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_33_711 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_700 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_744 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_733 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_722 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_777 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_766 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_33_755 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_32_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.DEC0.ABUF\[1\] A0BUF\[1\].X SLICE\[2\].RAM8.DEC0.A_buf\[1\] VDD VDD
+ VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_33_799 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfill_33_788 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0INV SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL0
+ SLICE\[0\].RAM8.WORD\[1\].W.BYTE\[3\].B.SEL0_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xtap_31_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_24_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WEBUF\[3\].__cell__ SLICE\[0\].RAM8.WEBUF\[3\].A SLICE\[3\].RAM8.WEBUF\[3\].X
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xtap_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.BIT\[7\].OBUF1 SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[0\].RAM8.WORD\[5\].W.BYTE\[1\].B.Q_WIRE\[7\] BYTE\[1\].FLOATBUF1\[15\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[0\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF1\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.BIT\[6\].genblk1.STORAGE DIBUF\[6\].X SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[6\].W.BYTE\[0\].B.Q_WIRE\[6\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.BIT\[7\].genblk1.STORAGE DIBUF\[15\].X SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.GCLK
+ SLICE\[0\].RAM8.WORD\[0\].W.BYTE\[1\].B.Q_WIRE\[7\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_26_43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XBYTE\[1\].FLOATBUF1\[8\].TE_BINV BYTE\[1\].FLOATBUF1\[10\].TE_B BYTE\[1\].FLOATBUF1\[8\].TE_BN
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_65 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_54 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[3\].OBUF1 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[3\] BYTE\[3\].FLOATBUF1\[27\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1INV SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[0\].B.SEL1_B VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
Xfill_26_98 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_26_87 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.BIT\[4\].OBUF0 SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.SEL0_B
+ SLICE\[2\].RAM8.WORD\[4\].W.BYTE\[1\].B.Q_WIRE\[4\] BYTE\[1\].FLOATBUF0\[12\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_9_106 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[1\].W.SEL1BUF SLICE\[2\].RAM8.WORD\[1\].W.SEL1 SLICE\[2\].RAM8.WORD\[1\].W.BYTE\[0\].B.SEL1
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfill_9_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_9_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_243 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_23_232 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.BIT\[1\].genblk1.STORAGE DIBUF\[25\].X SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[4\].W.BYTE\[3\].B.Q_WIRE\[1\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
XSLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.BIT\[0\].OBUF0 SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.SEL0_B
+ SLICE\[0\].RAM8.WORD\[7\].W.BYTE\[0\].B.Q_WIRE\[0\] BYTE\[0\].FLOATBUF0\[0\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
XSLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.BIT\[0\].genblk1.STORAGE DIBUF\[8\].X SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.GCLK
+ SLICE\[3\].RAM8.WORD\[2\].W.BYTE\[1\].B.Q_WIRE\[0\] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__latq_1
Xfill_0_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.BIT\[6\].OBUF0 SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.SEL0_B
+ SLICE\[1\].RAM8.WORD\[3\].W.BYTE\[3\].B.Q_WIRE\[6\] BYTE\[3\].FLOATBUF0\[30\].Z
+ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xfill_14_210 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_14_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_14_221 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtap_5_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XSLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.genblk1.CG SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.CLK_B
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.WE0_WIRE
+ SLICE\[3\].RAM8.WORD\[5\].W.BYTE\[0\].B.GCLK VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__icgtp_1
Xtap_5_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xtap_5_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfill_8_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_161 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_172 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_183 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfill_8_194 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XSLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.BIT\[0\].OBUF1 SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.SEL1_B
+ SLICE\[2\].RAM8.WORD\[3\].W.BYTE\[1\].B.Q_WIRE\[0\] BYTE\[1\].FLOATBUF1\[8\].Z VDD
+ VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__bufz_1
Xtap_10_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

